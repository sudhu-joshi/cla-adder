magic
tech scmos
timestamp 1732036114
<< nwell >>
rect -1 30 25 82
rect 31 30 57 82
rect 63 30 89 82
rect 95 30 121 82
rect 127 30 153 82
rect 161 30 187 82
<< ntransistor >>
rect 11 -100 13 0
rect 43 -106 45 -6
rect 75 -106 77 -6
rect 107 -106 109 -6
rect 139 -106 141 -6
rect 173 -39 175 1
<< ptransistor >>
rect 11 36 13 76
rect 43 36 45 76
rect 75 36 77 76
rect 107 36 109 76
rect 139 36 141 76
rect 173 36 175 76
<< ndiffusion >>
rect 10 -100 11 0
rect 13 -100 14 0
rect 42 -106 43 -6
rect 45 -106 46 -6
rect 74 -106 75 -6
rect 77 -106 78 -6
rect 106 -106 107 -6
rect 109 -106 110 -6
rect 138 -106 139 -6
rect 141 -106 142 -6
rect 172 -39 173 1
rect 175 -39 176 1
<< pdiffusion >>
rect 10 36 11 76
rect 13 36 14 76
rect 42 36 43 76
rect 45 36 46 76
rect 74 36 75 76
rect 77 36 78 76
rect 106 36 107 76
rect 109 36 110 76
rect 138 36 139 76
rect 141 36 142 76
rect 172 36 173 76
rect 175 36 176 76
<< ndcontact >>
rect 5 -100 10 0
rect 14 -100 19 0
rect 37 -106 42 -6
rect 46 -106 51 -6
rect 69 -106 74 -6
rect 78 -106 83 -6
rect 101 -106 106 -6
rect 110 -106 115 -6
rect 133 -106 138 -6
rect 142 -106 147 -6
rect 167 -39 172 1
rect 176 -39 181 1
<< pdcontact >>
rect 5 36 10 76
rect 14 36 19 76
rect 37 36 42 76
rect 46 36 51 76
rect 69 36 74 76
rect 78 36 83 76
rect 101 36 106 76
rect 110 36 115 76
rect 133 36 138 76
rect 142 36 147 76
rect 167 36 172 76
rect 176 36 181 76
<< polysilicon >>
rect 11 76 13 80
rect 43 76 45 80
rect 75 76 77 80
rect 107 76 109 80
rect 139 76 141 80
rect 173 76 175 80
rect 11 0 13 36
rect 43 22 45 36
rect 75 22 77 36
rect 107 22 109 36
rect 139 22 141 36
rect 43 -6 45 2
rect 75 -6 77 2
rect 107 -6 109 2
rect 139 -6 141 2
rect 173 1 175 36
rect 11 -103 13 -100
rect 173 -42 175 -39
rect 43 -110 45 -106
rect 75 -110 77 -106
rect 107 -110 109 -106
rect 139 -110 141 -106
<< polycontact >>
rect 6 22 11 27
rect 38 22 43 27
rect 70 22 75 27
rect 102 22 107 27
rect 134 22 139 27
rect 168 15 173 20
rect 38 -3 43 2
rect 70 -3 75 2
rect 102 -3 107 2
rect 134 -3 139 2
<< metal1 >>
rect -1 82 187 85
rect 5 76 10 82
rect 37 76 42 82
rect 69 76 74 82
rect 101 76 106 82
rect 133 76 138 82
rect 167 76 172 82
rect -1 22 6 27
rect 14 19 19 36
rect 35 22 38 27
rect 46 19 51 36
rect 67 22 70 27
rect 78 19 83 36
rect 99 22 102 27
rect 110 19 115 36
rect 131 22 134 27
rect 142 20 147 36
rect 176 22 181 36
rect 142 19 168 20
rect 14 16 168 19
rect 142 15 168 16
rect 176 17 187 22
rect 14 0 28 3
rect 5 -104 10 -100
rect 5 -110 19 -104
rect 24 -106 28 0
rect 35 -3 38 2
rect 46 -6 62 -2
rect 67 -3 70 2
rect 78 -6 94 -2
rect 99 -3 102 2
rect 110 -6 126 -2
rect 131 -3 134 2
rect 142 -6 147 15
rect 176 1 181 17
rect 58 -106 62 -6
rect 90 -106 94 -6
rect 24 -110 42 -106
rect 58 -110 74 -106
rect 90 -110 106 -106
rect 122 -107 126 -6
rect 167 -46 172 -39
rect 167 -50 181 -46
rect 133 -107 138 -106
rect 122 -110 138 -107
<< metal2 >>
rect 61 22 67 27
rect 61 17 64 22
rect -1 14 64 17
rect 61 2 64 14
rect 85 3 117 6
rect 61 -3 67 2
rect 85 1 88 3
rect 114 1 117 3
<< metal3 >>
rect 29 22 35 27
rect 29 21 32 22
rect -1 18 32 21
rect 29 2 32 18
rect 29 -3 35 2
<< metal4 >>
rect 96 13 99 27
rect -1 10 99 13
rect -1 3 85 6
rect 82 1 85 3
rect 96 -3 99 10
rect 128 6 131 27
rect 117 3 131 6
rect 117 1 120 3
rect 128 -3 131 3
<< metal5 >>
rect 96 13 99 27
rect -1 10 99 13
rect 96 -3 99 10
<< pad >>
rect 32 22 38 27
rect 64 22 70 27
rect 96 22 102 27
rect 128 22 134 27
rect 32 -3 38 2
rect 64 -3 70 2
rect 82 1 88 6
rect 96 -3 102 2
rect 114 1 120 6
rect 128 -3 134 2
<< labels >>
rlabel metal1 -1 22 6 27 3 a
rlabel metal3 -1 18 32 21 1 b
rlabel metal2 -1 14 64 17 1 c
rlabel metal5 -1 10 99 13 1 d
rlabel metal1 -1 82 187 85 5 vdd!
rlabel metal1 167 -50 172 -39 1 gnd!
rlabel metal1 176 1 181 36 1 out
rlabel metal1 5 -110 19 -104 1 gnd!
rlabel metal4 117 3 131 6 1 e
<< end >>
