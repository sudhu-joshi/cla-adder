.include TSMC_180nm.txt
.include subckt.txt

.param SUPPLY=1.8
.param LAMBDA = 0.09u
.param len = 2*LAMBDA
.param W_P = 20*LAMBDA
.param W_N = 10*LAMBDA

.global gnd vdd 
vdd vdd gnd 'SUPPLY'

* Input Pulses
VA A gnd pulse (0 SUPPLY 10ns .1ns .1ns 10ns 20ns)
VB B gnd pulse (0 SUPPLY 20ns .1ns .1ns 20ns 40ns)
* VC C gnd pulse (0 SUPPLY 40ns .1ns .1ns 40ns 80ns)
* VD D gnd pulse (0 SUPPLY 80ns .1ns .1ns 80ns 160ns)


* SPICE3 file created from or2.ext - technology: scmos

.option scale=0.09u

M1000 a_19_83# a vdd w_5_77# CMOSP w=60 l=2
+  ad=720 pd=264 as=720 ps=264
M1001 out a_19_15# vdd w_74_77# CMOSP w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1002 a_19_15# b gnd gnd CMOSN w=40 l=2
+  ad=480 pd=184 as=720 ps=276
M1003 a_19_15# b a_19_83# w_42_77# CMOSP w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1004 out a_19_15# gnd gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1005 a_19_15# a gnd gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_5_77# vdd 0.11fF
C1 gnd a_19_15# 0.89fF
C2 w_42_77# a_19_15# 0.09fF
C3 a_19_83# w_42_77# 0.11fF
C4 a_19_83# a_19_15# 0.65fF
C5 a_19_83# a 0.07fF
C6 a_19_83# w_5_77# 0.09fF
C7 w_74_77# vdd 0.11fF
C8 w_5_77# a 0.07fF
C9 out w_74_77# 0.09fF
C10 out vdd 0.65fF
C11 w_74_77# a_19_15# 0.07fF
C12 out gnd 0.41fF
C13 a_19_83# vdd 1.18fF
C14 out a_19_15# 0.07fF
C15 w_42_77# b 0.07fF
C16 a_19_15# b 0.05fF
C17 a_19_83# b 0.12fF
C18 a b 0.00fF
C19 gnd gnd 0.41fF
C20 out gnd 0.13fF
C21 a_19_83# gnd 0.42fF
C22 vdd gnd 0.27fF
C23 a_19_15# gnd 1.07fF
C24 b gnd 0.32fF
C25 a gnd 0.24fF
C26 w_74_77# gnd 0.12fF
C27 w_42_77# gnd 0.16fF
C28 w_5_77# gnd 0.16fF


* Simulation Setup
.tran 0.01ns 50ns
.control
    set hcopypscolor = 1
    set color0 = black
    set color1 = white
    run
    set curplottitle= o2_post
    plot v(A) v(B) v(out)+2

.endc
.end



