magic
tech scmos
timestamp 1733149062
<< nwell >>
rect -619 256 -593 308
rect -584 256 -558 308
rect -552 256 -526 308
rect -520 256 -494 308
rect -488 256 -462 308
rect -444 256 -418 308
rect -409 256 -383 308
rect -377 256 -351 308
rect -345 256 -319 308
rect -313 256 -287 308
rect -201 219 -149 245
rect -201 187 -149 213
rect -69 212 -17 238
rect -619 125 -593 177
rect -584 125 -558 177
rect -552 125 -526 177
rect -520 125 -494 177
rect -488 125 -462 177
rect -444 125 -418 177
rect -409 125 -383 177
rect -377 125 -351 177
rect -345 125 -319 177
rect -313 125 -287 177
rect -201 155 -149 181
rect -69 180 -17 206
rect 20 200 46 252
rect 52 200 78 252
rect 84 200 110 252
rect 131 225 157 277
rect 163 225 189 277
rect 195 225 221 277
rect 227 225 253 277
rect 458 192 484 403
rect 493 192 519 403
rect 528 192 554 403
rect 563 192 589 403
rect 598 192 624 403
rect -65 145 -13 171
rect 284 133 310 185
rect 316 133 342 185
rect 348 133 374 185
rect 380 133 406 185
rect 412 133 438 185
rect 630 183 656 235
rect 767 202 793 254
rect 802 202 828 254
rect 834 202 860 254
rect 866 202 892 254
rect 898 202 924 254
rect -201 91 -149 117
rect -201 59 -149 85
rect -69 84 -17 110
rect -619 -7 -593 45
rect -584 -7 -558 45
rect -552 -7 -526 45
rect -520 -7 -494 45
rect -488 -7 -462 45
rect -444 -7 -418 45
rect -409 -7 -383 45
rect -377 -7 -351 45
rect -345 -7 -319 45
rect -313 -7 -287 45
rect -201 27 -149 53
rect -69 52 -17 78
rect 28 52 54 104
rect 60 52 86 104
rect 92 52 118 104
rect 134 68 160 120
rect 166 68 192 120
rect 198 68 224 120
rect 230 68 256 120
rect 662 109 688 161
rect 694 109 720 161
rect 729 113 755 165
rect 445 45 471 97
rect 477 45 503 97
rect 509 45 535 97
rect 541 45 567 97
rect 573 45 599 97
rect 607 45 633 97
rect 767 70 793 122
rect 802 70 828 122
rect 834 70 860 122
rect 866 70 892 122
rect 898 70 924 122
rect -65 17 -13 43
rect -201 -37 -149 -11
rect -201 -69 -149 -43
rect -69 -44 -17 -18
rect -619 -138 -593 -86
rect -584 -138 -558 -86
rect -552 -138 -526 -86
rect -520 -138 -494 -86
rect -488 -138 -462 -86
rect -444 -138 -418 -86
rect -409 -138 -383 -86
rect -377 -138 -351 -86
rect -345 -138 -319 -86
rect -313 -138 -287 -86
rect -201 -101 -149 -75
rect -69 -76 -17 -50
rect -65 -111 -13 -85
rect 30 -94 56 -42
rect 62 -94 88 -42
rect 94 -94 120 -42
rect 126 -94 152 -42
rect 276 -55 302 -3
rect 308 -55 334 -3
rect 340 -55 366 -3
rect 372 -55 398 -3
rect 404 -55 430 -3
rect 662 -36 688 16
rect 694 -36 720 16
rect 729 -32 755 20
rect 162 -110 188 -58
rect 194 -110 220 -58
rect 226 -110 252 -58
rect 767 -61 793 -9
rect 802 -61 828 -9
rect 834 -61 860 -9
rect 866 -61 892 -9
rect 898 -61 924 -9
rect -201 -165 -149 -139
rect -201 -197 -149 -171
rect -69 -172 -17 -146
rect -201 -229 -149 -203
rect -69 -204 -17 -178
rect -65 -239 -13 -213
rect 30 -247 56 -195
rect 62 -247 88 -195
rect 94 -247 120 -195
rect 126 -258 152 -206
rect 163 -258 189 -206
rect 195 -258 221 -206
rect 265 -249 291 -177
rect 300 -249 326 -177
rect 335 -249 361 -177
rect 367 -256 393 -204
rect 427 -235 453 -143
rect 462 -235 488 -143
rect 497 -235 523 -143
rect 532 -235 558 -143
rect 639 -183 665 -131
rect 671 -183 697 -131
rect 706 -179 732 -127
rect 564 -242 590 -190
rect 767 -193 793 -141
rect 802 -193 828 -141
rect 834 -193 860 -141
rect 866 -193 892 -141
rect 898 -193 924 -141
rect -183 -322 -157 -270
rect -148 -322 -122 -270
rect -116 -322 -90 -270
rect -84 -322 -58 -270
rect -52 -322 -26 -270
rect 639 -328 665 -276
rect 671 -328 697 -276
rect 706 -324 732 -272
rect 767 -324 793 -272
rect 802 -324 828 -272
rect 834 -324 860 -272
rect 866 -324 892 -272
rect 898 -324 924 -272
<< ntransistor >>
rect -607 206 -605 236
rect -589 202 -587 232
rect -566 202 -564 232
rect -536 202 -534 232
rect -513 202 -511 232
rect -476 212 -474 242
rect -432 206 -430 236
rect -414 202 -412 232
rect -391 202 -389 232
rect -361 202 -359 232
rect -338 202 -336 232
rect -301 212 -299 242
rect -263 231 -223 233
rect -130 224 -90 226
rect -266 199 -226 201
rect -130 192 -90 194
rect -262 167 -222 169
rect -130 157 -90 159
rect 32 138 34 178
rect 64 135 66 175
rect 96 139 98 179
rect 143 143 145 203
rect 175 137 177 197
rect 207 137 209 197
rect 239 164 241 204
rect -607 75 -605 105
rect -589 71 -587 101
rect -566 71 -564 101
rect -536 71 -534 101
rect -513 71 -511 101
rect -476 81 -474 111
rect -432 75 -430 105
rect -414 71 -412 101
rect -391 71 -389 101
rect -361 71 -359 101
rect -338 71 -336 101
rect -301 81 -299 111
rect -263 103 -223 105
rect -130 96 -90 98
rect -266 71 -226 73
rect -130 64 -90 66
rect -262 39 -222 41
rect -130 29 -90 31
rect -607 -57 -605 -27
rect -589 -61 -587 -31
rect -566 -61 -564 -31
rect -536 -61 -534 -31
rect -513 -61 -511 -31
rect -476 -51 -474 -21
rect 40 -10 42 30
rect 72 -13 74 27
rect 104 -9 106 31
rect 146 -14 148 46
rect -432 -57 -430 -27
rect -414 -61 -412 -31
rect -391 -61 -389 -31
rect -361 -61 -359 -31
rect -338 -61 -336 -31
rect -301 -51 -299 -21
rect 178 -20 180 40
rect 210 -20 212 40
rect 242 7 244 47
rect 296 29 298 109
rect 470 117 472 157
rect 505 116 507 156
rect 540 116 542 156
rect 575 116 577 156
rect 610 116 612 156
rect 642 116 644 156
rect 779 152 781 182
rect 797 148 799 178
rect 820 148 822 178
rect 850 148 852 178
rect 873 148 875 178
rect 910 158 912 188
rect 328 23 330 103
rect 360 23 362 103
rect 392 23 394 103
rect 424 70 426 110
rect -263 -25 -223 -23
rect -130 -32 -90 -30
rect -266 -57 -226 -55
rect -130 -64 -90 -62
rect -262 -89 -222 -87
rect -130 -99 -90 -97
rect -607 -188 -605 -158
rect -589 -192 -587 -162
rect -566 -192 -564 -162
rect -536 -192 -534 -162
rect -513 -192 -511 -162
rect -476 -182 -474 -152
rect -432 -188 -430 -158
rect -414 -192 -412 -162
rect -391 -192 -389 -162
rect -361 -192 -359 -162
rect -338 -192 -336 -162
rect -301 -182 -299 -152
rect -263 -153 -223 -151
rect -130 -160 -90 -158
rect 42 -176 44 -116
rect 74 -182 76 -122
rect 106 -182 108 -122
rect 138 -155 140 -115
rect 174 -172 176 -132
rect 206 -175 208 -135
rect 238 -171 240 -131
rect 288 -159 290 -79
rect 320 -165 322 -85
rect 352 -165 354 -85
rect 384 -165 386 -85
rect 416 -118 418 -78
rect 457 -85 459 15
rect 674 48 676 88
rect 706 48 708 88
rect 741 48 743 88
rect 779 20 781 50
rect 489 -91 491 9
rect 521 -91 523 9
rect 553 -91 555 9
rect 585 -91 587 9
rect 619 -24 621 16
rect 797 16 799 46
rect 820 16 822 46
rect 850 16 852 46
rect 873 16 875 46
rect 910 26 912 56
rect 674 -97 676 -57
rect 706 -97 708 -57
rect 741 -97 743 -57
rect 779 -111 781 -81
rect 797 -115 799 -85
rect 820 -115 822 -85
rect 850 -115 852 -85
rect 873 -115 875 -85
rect 910 -105 912 -75
rect -266 -185 -226 -183
rect -130 -192 -90 -190
rect -262 -217 -222 -215
rect -130 -227 -90 -225
rect 42 -309 44 -269
rect 74 -312 76 -272
rect 106 -308 108 -268
rect 138 -320 140 -280
rect 175 -320 177 -280
rect 207 -319 209 -279
rect 277 -316 279 -276
rect 312 -317 314 -277
rect 347 -317 349 -277
rect 379 -317 381 -277
rect 439 -306 441 -266
rect 651 -244 653 -204
rect 683 -244 685 -204
rect 718 -244 720 -204
rect 779 -243 781 -213
rect 797 -247 799 -217
rect 820 -247 822 -217
rect 850 -247 852 -217
rect 873 -247 875 -217
rect 910 -237 912 -207
rect 474 -307 476 -267
rect 509 -307 511 -267
rect 544 -307 546 -267
rect 576 -307 578 -267
rect -171 -372 -169 -342
rect -153 -376 -151 -346
rect -130 -376 -128 -346
rect -100 -376 -98 -346
rect -77 -376 -75 -346
rect -40 -366 -38 -336
rect 651 -389 653 -349
rect 683 -389 685 -349
rect 718 -389 720 -349
rect 779 -374 781 -344
rect 797 -378 799 -348
rect 820 -378 822 -348
rect 850 -378 852 -348
rect 873 -378 875 -348
rect 910 -368 912 -338
<< ptransistor >>
rect -607 262 -605 302
rect -572 262 -570 302
rect -540 262 -538 302
rect -508 262 -506 302
rect -476 262 -474 302
rect -432 262 -430 302
rect -397 262 -395 302
rect -365 262 -363 302
rect -333 262 -331 302
rect -301 262 -299 302
rect -195 231 -155 233
rect -63 224 -23 226
rect 32 206 34 246
rect 64 206 66 246
rect 96 206 98 246
rect 143 231 145 271
rect 175 231 177 271
rect 207 231 209 271
rect 239 231 241 271
rect -195 199 -155 201
rect -63 192 -23 194
rect -607 131 -605 171
rect -572 131 -570 171
rect -540 131 -538 171
rect -508 131 -506 171
rect -476 131 -474 171
rect -432 131 -430 171
rect -397 131 -395 171
rect -365 131 -363 171
rect -333 131 -331 171
rect -301 131 -299 171
rect -195 167 -155 169
rect -59 157 -19 159
rect 470 198 472 397
rect 505 198 507 397
rect 540 198 542 397
rect 575 198 577 397
rect 610 198 612 397
rect 296 139 298 179
rect 328 139 330 179
rect 360 139 362 179
rect 392 139 394 179
rect 424 139 426 179
rect 642 189 644 229
rect 779 208 781 248
rect 814 208 816 248
rect 846 208 848 248
rect 878 208 880 248
rect 910 208 912 248
rect -195 103 -155 105
rect -63 96 -23 98
rect -195 71 -155 73
rect -63 64 -23 66
rect 40 58 42 98
rect 72 58 74 98
rect 104 58 106 98
rect 146 74 148 114
rect 178 74 180 114
rect 210 74 212 114
rect 242 74 244 114
rect -195 39 -155 41
rect -607 -1 -605 39
rect -572 -1 -570 39
rect -540 -1 -538 39
rect -508 -1 -506 39
rect -476 -1 -474 39
rect -432 -1 -430 39
rect -397 -1 -395 39
rect -365 -1 -363 39
rect -333 -1 -331 39
rect -301 -1 -299 39
rect -59 29 -19 31
rect 674 115 676 155
rect 706 115 708 155
rect 741 119 743 159
rect 457 51 459 91
rect 489 51 491 91
rect 521 51 523 91
rect 553 51 555 91
rect 585 51 587 91
rect 619 51 621 91
rect -195 -25 -155 -23
rect -63 -32 -23 -30
rect -195 -57 -155 -55
rect -63 -64 -23 -62
rect -195 -89 -155 -87
rect 42 -88 44 -48
rect 74 -88 76 -48
rect 106 -88 108 -48
rect 138 -88 140 -48
rect 288 -49 290 -9
rect 320 -49 322 -9
rect 352 -49 354 -9
rect 384 -49 386 -9
rect 416 -49 418 -9
rect -607 -132 -605 -92
rect -572 -132 -570 -92
rect -540 -132 -538 -92
rect -508 -132 -506 -92
rect -476 -132 -474 -92
rect -432 -132 -430 -92
rect -397 -132 -395 -92
rect -365 -132 -363 -92
rect -333 -132 -331 -92
rect -301 -132 -299 -92
rect -59 -99 -19 -97
rect -195 -153 -155 -151
rect -63 -160 -23 -158
rect 174 -104 176 -64
rect 206 -104 208 -64
rect 238 -104 240 -64
rect 779 76 781 116
rect 814 76 816 116
rect 846 76 848 116
rect 878 76 880 116
rect 910 76 912 116
rect 674 -30 676 10
rect 706 -30 708 10
rect 741 -26 743 14
rect 779 -55 781 -15
rect 814 -55 816 -15
rect 846 -55 848 -15
rect 878 -55 880 -15
rect 910 -55 912 -15
rect -195 -185 -155 -183
rect -63 -192 -23 -190
rect -195 -217 -155 -215
rect -59 -227 -19 -225
rect 42 -241 44 -201
rect 74 -241 76 -201
rect 106 -241 108 -201
rect -171 -316 -169 -276
rect -136 -316 -134 -276
rect -104 -316 -102 -276
rect -72 -316 -70 -276
rect -40 -316 -38 -276
rect 138 -252 140 -212
rect 175 -252 177 -212
rect 207 -252 209 -212
rect 277 -243 279 -183
rect 312 -243 314 -183
rect 347 -243 349 -183
rect 379 -250 381 -210
rect 439 -229 441 -149
rect 474 -229 476 -149
rect 509 -229 511 -149
rect 544 -229 546 -149
rect 651 -177 653 -137
rect 683 -177 685 -137
rect 718 -173 720 -133
rect 576 -236 578 -196
rect 779 -187 781 -147
rect 814 -187 816 -147
rect 846 -187 848 -147
rect 878 -187 880 -147
rect 910 -187 912 -147
rect 651 -322 653 -282
rect 683 -322 685 -282
rect 718 -318 720 -278
rect 779 -318 781 -278
rect 814 -318 816 -278
rect 846 -318 848 -278
rect 878 -318 880 -278
rect 910 -318 912 -278
<< ndiffusion >>
rect -608 206 -607 236
rect -605 206 -604 236
rect -590 202 -589 232
rect -587 202 -586 232
rect -567 202 -566 232
rect -564 202 -563 232
rect -537 202 -536 232
rect -534 202 -533 232
rect -514 202 -513 232
rect -511 202 -510 232
rect -477 212 -476 242
rect -474 212 -473 242
rect -433 206 -432 236
rect -430 206 -429 236
rect -415 202 -414 232
rect -412 202 -411 232
rect -392 202 -391 232
rect -389 202 -388 232
rect -362 202 -361 232
rect -359 202 -358 232
rect -339 202 -338 232
rect -336 202 -335 232
rect -302 212 -301 242
rect -299 212 -298 242
rect -263 233 -223 234
rect -263 230 -223 231
rect -130 226 -90 227
rect -130 223 -90 224
rect -266 201 -226 202
rect -266 198 -226 199
rect -130 194 -90 195
rect -130 191 -90 192
rect -262 169 -222 170
rect -262 166 -222 167
rect -130 159 -90 160
rect -130 156 -90 157
rect 31 138 32 178
rect 34 138 35 178
rect 63 135 64 175
rect 66 135 67 175
rect 95 139 96 179
rect 98 139 99 179
rect 142 143 143 203
rect 145 143 146 203
rect 174 137 175 197
rect 177 137 178 197
rect 206 137 207 197
rect 209 137 210 197
rect 238 164 239 204
rect 241 164 242 204
rect -608 75 -607 105
rect -605 75 -604 105
rect -590 71 -589 101
rect -587 71 -586 101
rect -567 71 -566 101
rect -564 71 -563 101
rect -537 71 -536 101
rect -534 71 -533 101
rect -514 71 -513 101
rect -511 71 -510 101
rect -477 81 -476 111
rect -474 81 -473 111
rect -433 75 -432 105
rect -430 75 -429 105
rect -415 71 -414 101
rect -412 71 -411 101
rect -392 71 -391 101
rect -389 71 -388 101
rect -362 71 -361 101
rect -359 71 -358 101
rect -339 71 -338 101
rect -336 71 -335 101
rect -302 81 -301 111
rect -299 81 -298 111
rect -263 105 -223 106
rect -263 102 -223 103
rect -130 98 -90 99
rect -130 95 -90 96
rect -266 73 -226 74
rect -266 70 -226 71
rect -130 66 -90 67
rect -130 63 -90 64
rect -262 41 -222 42
rect -262 38 -222 39
rect -130 31 -90 32
rect -130 28 -90 29
rect -608 -57 -607 -27
rect -605 -57 -604 -27
rect -590 -61 -589 -31
rect -587 -61 -586 -31
rect -567 -61 -566 -31
rect -564 -61 -563 -31
rect -537 -61 -536 -31
rect -534 -61 -533 -31
rect -514 -61 -513 -31
rect -511 -61 -510 -31
rect -477 -51 -476 -21
rect -474 -51 -473 -21
rect 39 -10 40 30
rect 42 -10 43 30
rect 71 -13 72 27
rect 74 -13 75 27
rect 103 -9 104 31
rect 106 -9 107 31
rect 145 -14 146 46
rect 148 -14 149 46
rect -433 -57 -432 -27
rect -430 -57 -429 -27
rect -415 -61 -414 -31
rect -412 -61 -411 -31
rect -392 -61 -391 -31
rect -389 -61 -388 -31
rect -362 -61 -361 -31
rect -359 -61 -358 -31
rect -339 -61 -338 -31
rect -336 -61 -335 -31
rect -302 -51 -301 -21
rect -299 -51 -298 -21
rect -263 -23 -223 -22
rect 177 -20 178 40
rect 180 -20 181 40
rect 209 -20 210 40
rect 212 -20 213 40
rect 241 7 242 47
rect 244 7 245 47
rect 295 29 296 109
rect 298 29 299 109
rect 469 117 470 157
rect 472 117 473 157
rect 504 116 505 156
rect 507 116 508 156
rect 539 116 540 156
rect 542 116 543 156
rect 574 116 575 156
rect 577 116 578 156
rect 609 116 610 156
rect 612 116 613 156
rect 641 116 642 156
rect 644 116 645 156
rect 778 152 779 182
rect 781 152 782 182
rect 796 148 797 178
rect 799 148 800 178
rect 819 148 820 178
rect 822 148 823 178
rect 849 148 850 178
rect 852 148 853 178
rect 872 148 873 178
rect 875 148 876 178
rect 909 158 910 188
rect 912 158 913 188
rect 327 23 328 103
rect 330 23 331 103
rect 359 23 360 103
rect 362 23 363 103
rect 391 23 392 103
rect 394 23 395 103
rect 423 70 424 110
rect 426 70 427 110
rect -263 -26 -223 -25
rect -130 -30 -90 -29
rect -130 -33 -90 -32
rect -266 -55 -226 -54
rect -266 -58 -226 -57
rect -130 -62 -90 -61
rect -130 -65 -90 -64
rect -262 -87 -222 -86
rect -262 -90 -222 -89
rect -130 -97 -90 -96
rect -130 -100 -90 -99
rect -608 -188 -607 -158
rect -605 -188 -604 -158
rect -590 -192 -589 -162
rect -587 -192 -586 -162
rect -567 -192 -566 -162
rect -564 -192 -563 -162
rect -537 -192 -536 -162
rect -534 -192 -533 -162
rect -514 -192 -513 -162
rect -511 -192 -510 -162
rect -477 -182 -476 -152
rect -474 -182 -473 -152
rect -263 -151 -223 -150
rect -433 -188 -432 -158
rect -430 -188 -429 -158
rect -415 -192 -414 -162
rect -412 -192 -411 -162
rect -392 -192 -391 -162
rect -389 -192 -388 -162
rect -362 -192 -361 -162
rect -359 -192 -358 -162
rect -339 -192 -338 -162
rect -336 -192 -335 -162
rect -302 -182 -301 -152
rect -299 -182 -298 -152
rect -263 -154 -223 -153
rect -130 -158 -90 -157
rect -130 -161 -90 -160
rect 41 -176 42 -116
rect 44 -176 45 -116
rect -266 -183 -226 -182
rect 73 -182 74 -122
rect 76 -182 77 -122
rect 105 -182 106 -122
rect 108 -182 109 -122
rect 137 -155 138 -115
rect 140 -155 141 -115
rect 173 -172 174 -132
rect 176 -172 177 -132
rect 205 -175 206 -135
rect 208 -175 209 -135
rect 237 -171 238 -131
rect 240 -171 241 -131
rect 287 -159 288 -79
rect 290 -159 291 -79
rect 319 -165 320 -85
rect 322 -165 323 -85
rect 351 -165 352 -85
rect 354 -165 355 -85
rect 383 -165 384 -85
rect 386 -165 387 -85
rect 415 -118 416 -78
rect 418 -118 419 -78
rect 456 -85 457 15
rect 459 -85 460 15
rect 673 48 674 88
rect 676 48 677 88
rect 705 48 706 88
rect 708 48 709 88
rect 740 48 741 88
rect 743 48 744 88
rect 778 20 779 50
rect 781 20 782 50
rect 488 -91 489 9
rect 491 -91 492 9
rect 520 -91 521 9
rect 523 -91 524 9
rect 552 -91 553 9
rect 555 -91 556 9
rect 584 -91 585 9
rect 587 -91 588 9
rect 618 -24 619 16
rect 621 -24 622 16
rect 796 16 797 46
rect 799 16 800 46
rect 819 16 820 46
rect 822 16 823 46
rect 849 16 850 46
rect 852 16 853 46
rect 872 16 873 46
rect 875 16 876 46
rect 909 26 910 56
rect 912 26 913 56
rect 673 -97 674 -57
rect 676 -97 677 -57
rect 705 -97 706 -57
rect 708 -97 709 -57
rect 740 -97 741 -57
rect 743 -97 744 -57
rect 778 -111 779 -81
rect 781 -111 782 -81
rect 796 -115 797 -85
rect 799 -115 800 -85
rect 819 -115 820 -85
rect 822 -115 823 -85
rect 849 -115 850 -85
rect 852 -115 853 -85
rect 872 -115 873 -85
rect 875 -115 876 -85
rect 909 -105 910 -75
rect 912 -105 913 -75
rect -266 -186 -226 -185
rect -130 -190 -90 -189
rect -130 -193 -90 -192
rect -262 -215 -222 -214
rect -262 -218 -222 -217
rect -130 -225 -90 -224
rect -130 -228 -90 -227
rect 41 -309 42 -269
rect 44 -309 45 -269
rect 73 -312 74 -272
rect 76 -312 77 -272
rect 105 -308 106 -268
rect 108 -308 109 -268
rect 137 -320 138 -280
rect 140 -320 141 -280
rect 174 -320 175 -280
rect 177 -320 178 -280
rect 206 -319 207 -279
rect 209 -319 210 -279
rect 276 -316 277 -276
rect 279 -316 280 -276
rect 311 -317 312 -277
rect 314 -317 315 -277
rect 346 -317 347 -277
rect 349 -317 350 -277
rect 378 -317 379 -277
rect 381 -317 382 -277
rect 438 -306 439 -266
rect 441 -306 442 -266
rect 650 -244 651 -204
rect 653 -244 654 -204
rect 682 -244 683 -204
rect 685 -244 686 -204
rect 717 -244 718 -204
rect 720 -244 721 -204
rect 778 -243 779 -213
rect 781 -243 782 -213
rect 796 -247 797 -217
rect 799 -247 800 -217
rect 819 -247 820 -217
rect 822 -247 823 -217
rect 849 -247 850 -217
rect 852 -247 853 -217
rect 872 -247 873 -217
rect 875 -247 876 -217
rect 909 -237 910 -207
rect 912 -237 913 -207
rect 473 -307 474 -267
rect 476 -307 477 -267
rect 508 -307 509 -267
rect 511 -307 512 -267
rect 543 -307 544 -267
rect 546 -307 547 -267
rect 575 -307 576 -267
rect 578 -307 579 -267
rect -172 -372 -171 -342
rect -169 -372 -168 -342
rect -154 -376 -153 -346
rect -151 -376 -150 -346
rect -131 -376 -130 -346
rect -128 -376 -127 -346
rect -101 -376 -100 -346
rect -98 -376 -97 -346
rect -78 -376 -77 -346
rect -75 -376 -74 -346
rect -41 -366 -40 -336
rect -38 -366 -37 -336
rect 650 -389 651 -349
rect 653 -389 654 -349
rect 682 -389 683 -349
rect 685 -389 686 -349
rect 717 -389 718 -349
rect 720 -389 721 -349
rect 778 -374 779 -344
rect 781 -374 782 -344
rect 796 -378 797 -348
rect 799 -378 800 -348
rect 819 -378 820 -348
rect 822 -378 823 -348
rect 849 -378 850 -348
rect 852 -378 853 -348
rect 872 -378 873 -348
rect 875 -378 876 -348
rect 909 -368 910 -338
rect 912 -368 913 -338
<< pdiffusion >>
rect -608 262 -607 302
rect -605 262 -604 302
rect -573 262 -572 302
rect -570 262 -569 302
rect -541 262 -540 302
rect -538 262 -537 302
rect -509 262 -508 302
rect -506 262 -505 302
rect -477 262 -476 302
rect -474 262 -473 302
rect -433 262 -432 302
rect -430 262 -429 302
rect -398 262 -397 302
rect -395 262 -394 302
rect -366 262 -365 302
rect -363 262 -362 302
rect -334 262 -333 302
rect -331 262 -330 302
rect -302 262 -301 302
rect -299 262 -298 302
rect -195 233 -155 234
rect -195 230 -155 231
rect -63 226 -23 227
rect -63 223 -23 224
rect 31 206 32 246
rect 34 206 35 246
rect 63 206 64 246
rect 66 206 67 246
rect 95 206 96 246
rect 98 206 99 246
rect 142 231 143 271
rect 145 231 146 271
rect 174 231 175 271
rect 177 231 178 271
rect 206 231 207 271
rect 209 231 210 271
rect 238 231 239 271
rect 241 231 242 271
rect -195 201 -155 202
rect -195 198 -155 199
rect -63 194 -23 195
rect -63 191 -23 192
rect -608 131 -607 171
rect -605 131 -604 171
rect -573 131 -572 171
rect -570 131 -569 171
rect -541 131 -540 171
rect -538 131 -537 171
rect -509 131 -508 171
rect -506 131 -505 171
rect -477 131 -476 171
rect -474 131 -473 171
rect -433 131 -432 171
rect -430 131 -429 171
rect -398 131 -397 171
rect -395 131 -394 171
rect -366 131 -365 171
rect -363 131 -362 171
rect -334 131 -333 171
rect -331 131 -330 171
rect -302 131 -301 171
rect -299 131 -298 171
rect -195 169 -155 170
rect -195 166 -155 167
rect -59 159 -19 160
rect -59 156 -19 157
rect 469 198 470 397
rect 472 198 473 397
rect 504 198 505 397
rect 507 198 508 397
rect 539 198 540 397
rect 542 198 543 397
rect 574 198 575 397
rect 577 198 578 397
rect 609 198 610 397
rect 612 198 613 397
rect 295 139 296 179
rect 298 139 299 179
rect 327 139 328 179
rect 330 139 331 179
rect 359 139 360 179
rect 362 139 363 179
rect 391 139 392 179
rect 394 139 395 179
rect 423 139 424 179
rect 426 139 427 179
rect 641 189 642 229
rect 644 189 645 229
rect 778 208 779 248
rect 781 208 782 248
rect 813 208 814 248
rect 816 208 817 248
rect 845 208 846 248
rect 848 208 849 248
rect 877 208 878 248
rect 880 208 881 248
rect 909 208 910 248
rect 912 208 913 248
rect -195 105 -155 106
rect -195 102 -155 103
rect -63 98 -23 99
rect -63 95 -23 96
rect -195 73 -155 74
rect -195 70 -155 71
rect -63 66 -23 67
rect -63 63 -23 64
rect 39 58 40 98
rect 42 58 43 98
rect 71 58 72 98
rect 74 58 75 98
rect 103 58 104 98
rect 106 58 107 98
rect 145 74 146 114
rect 148 74 149 114
rect 177 74 178 114
rect 180 74 181 114
rect 209 74 210 114
rect 212 74 213 114
rect 241 74 242 114
rect 244 74 245 114
rect -195 41 -155 42
rect -608 -1 -607 39
rect -605 -1 -604 39
rect -573 -1 -572 39
rect -570 -1 -569 39
rect -541 -1 -540 39
rect -538 -1 -537 39
rect -509 -1 -508 39
rect -506 -1 -505 39
rect -477 -1 -476 39
rect -474 -1 -473 39
rect -433 -1 -432 39
rect -430 -1 -429 39
rect -398 -1 -397 39
rect -395 -1 -394 39
rect -366 -1 -365 39
rect -363 -1 -362 39
rect -334 -1 -333 39
rect -331 -1 -330 39
rect -302 -1 -301 39
rect -299 -1 -298 39
rect -195 38 -155 39
rect -59 31 -19 32
rect -59 28 -19 29
rect 673 115 674 155
rect 676 115 677 155
rect 705 115 706 155
rect 708 115 709 155
rect 740 119 741 159
rect 743 119 744 159
rect 456 51 457 91
rect 459 51 460 91
rect 488 51 489 91
rect 491 51 492 91
rect 520 51 521 91
rect 523 51 524 91
rect 552 51 553 91
rect 555 51 556 91
rect 584 51 585 91
rect 587 51 588 91
rect 618 51 619 91
rect 621 51 622 91
rect -195 -23 -155 -22
rect -195 -26 -155 -25
rect -63 -30 -23 -29
rect -63 -33 -23 -32
rect -195 -55 -155 -54
rect -195 -58 -155 -57
rect -63 -62 -23 -61
rect -63 -65 -23 -64
rect -195 -87 -155 -86
rect 41 -88 42 -48
rect 44 -88 45 -48
rect 73 -88 74 -48
rect 76 -88 77 -48
rect 105 -88 106 -48
rect 108 -88 109 -48
rect 137 -88 138 -48
rect 140 -88 141 -48
rect 287 -49 288 -9
rect 290 -49 291 -9
rect 319 -49 320 -9
rect 322 -49 323 -9
rect 351 -49 352 -9
rect 354 -49 355 -9
rect 383 -49 384 -9
rect 386 -49 387 -9
rect 415 -49 416 -9
rect 418 -49 419 -9
rect -608 -132 -607 -92
rect -605 -132 -604 -92
rect -573 -132 -572 -92
rect -570 -132 -569 -92
rect -541 -132 -540 -92
rect -538 -132 -537 -92
rect -509 -132 -508 -92
rect -506 -132 -505 -92
rect -477 -132 -476 -92
rect -474 -132 -473 -92
rect -433 -132 -432 -92
rect -430 -132 -429 -92
rect -398 -132 -397 -92
rect -395 -132 -394 -92
rect -366 -132 -365 -92
rect -363 -132 -362 -92
rect -334 -132 -333 -92
rect -331 -132 -330 -92
rect -302 -132 -301 -92
rect -299 -132 -298 -92
rect -195 -90 -155 -89
rect -59 -97 -19 -96
rect -59 -100 -19 -99
rect -195 -151 -155 -150
rect -195 -154 -155 -153
rect -63 -158 -23 -157
rect -63 -161 -23 -160
rect 173 -104 174 -64
rect 176 -104 177 -64
rect 205 -104 206 -64
rect 208 -104 209 -64
rect 237 -104 238 -64
rect 240 -104 241 -64
rect 778 76 779 116
rect 781 76 782 116
rect 813 76 814 116
rect 816 76 817 116
rect 845 76 846 116
rect 848 76 849 116
rect 877 76 878 116
rect 880 76 881 116
rect 909 76 910 116
rect 912 76 913 116
rect 673 -30 674 10
rect 676 -30 677 10
rect 705 -30 706 10
rect 708 -30 709 10
rect 740 -26 741 14
rect 743 -26 744 14
rect 778 -55 779 -15
rect 781 -55 782 -15
rect 813 -55 814 -15
rect 816 -55 817 -15
rect 845 -55 846 -15
rect 848 -55 849 -15
rect 877 -55 878 -15
rect 880 -55 881 -15
rect 909 -55 910 -15
rect 912 -55 913 -15
rect -195 -183 -155 -182
rect -195 -186 -155 -185
rect -63 -190 -23 -189
rect -63 -193 -23 -192
rect -195 -215 -155 -214
rect -195 -218 -155 -217
rect -59 -225 -19 -224
rect -59 -228 -19 -227
rect 41 -241 42 -201
rect 44 -241 45 -201
rect 73 -241 74 -201
rect 76 -241 77 -201
rect 105 -241 106 -201
rect 108 -241 109 -201
rect -172 -316 -171 -276
rect -169 -316 -168 -276
rect -137 -316 -136 -276
rect -134 -316 -133 -276
rect -105 -316 -104 -276
rect -102 -316 -101 -276
rect -73 -316 -72 -276
rect -70 -316 -69 -276
rect -41 -316 -40 -276
rect -38 -316 -37 -276
rect 137 -252 138 -212
rect 140 -252 141 -212
rect 174 -252 175 -212
rect 177 -252 178 -212
rect 206 -252 207 -212
rect 209 -252 210 -212
rect 276 -243 277 -183
rect 279 -243 280 -183
rect 311 -243 312 -183
rect 314 -243 315 -183
rect 346 -243 347 -183
rect 349 -243 350 -183
rect 378 -250 379 -210
rect 381 -250 382 -210
rect 438 -229 439 -149
rect 441 -229 442 -149
rect 473 -229 474 -149
rect 476 -229 477 -149
rect 508 -229 509 -149
rect 511 -229 512 -149
rect 543 -229 544 -149
rect 546 -229 547 -149
rect 650 -177 651 -137
rect 653 -177 654 -137
rect 682 -177 683 -137
rect 685 -177 686 -137
rect 717 -173 718 -133
rect 720 -173 721 -133
rect 575 -236 576 -196
rect 578 -236 579 -196
rect 778 -187 779 -147
rect 781 -187 782 -147
rect 813 -187 814 -147
rect 816 -187 817 -147
rect 845 -187 846 -147
rect 848 -187 849 -147
rect 877 -187 878 -147
rect 880 -187 881 -147
rect 909 -187 910 -147
rect 912 -187 913 -147
rect 650 -322 651 -282
rect 653 -322 654 -282
rect 682 -322 683 -282
rect 685 -322 686 -282
rect 717 -318 718 -278
rect 720 -318 721 -278
rect 778 -318 779 -278
rect 781 -318 782 -278
rect 813 -318 814 -278
rect 816 -318 817 -278
rect 845 -318 846 -278
rect 848 -318 849 -278
rect 877 -318 878 -278
rect 880 -318 881 -278
rect 909 -318 910 -278
rect 912 -318 913 -278
<< ndcontact >>
rect -613 206 -608 236
rect -604 206 -599 236
rect -595 202 -590 232
rect -586 202 -581 232
rect -572 202 -567 232
rect -563 202 -558 232
rect -542 202 -537 232
rect -533 202 -528 232
rect -519 202 -514 232
rect -510 202 -505 232
rect -482 212 -477 242
rect -473 212 -468 242
rect -438 206 -433 236
rect -429 206 -424 236
rect -420 202 -415 232
rect -411 202 -406 232
rect -397 202 -392 232
rect -388 202 -383 232
rect -367 202 -362 232
rect -358 202 -353 232
rect -344 202 -339 232
rect -335 202 -330 232
rect -307 212 -302 242
rect -298 212 -293 242
rect -263 234 -223 239
rect -263 225 -223 230
rect -130 227 -90 232
rect -130 218 -90 223
rect -266 202 -226 207
rect -266 193 -226 198
rect -130 195 -90 200
rect -130 186 -90 191
rect -262 170 -222 175
rect -262 161 -222 166
rect -130 160 -90 165
rect -130 151 -90 156
rect 26 138 31 178
rect 35 138 40 178
rect 58 135 63 175
rect 67 135 72 175
rect 90 139 95 179
rect 99 139 104 179
rect 137 143 142 203
rect 146 143 151 203
rect 169 137 174 197
rect 178 137 183 197
rect 201 137 206 197
rect 210 137 215 197
rect 233 164 238 204
rect 242 164 247 204
rect -613 75 -608 105
rect -604 75 -599 105
rect -595 71 -590 101
rect -586 71 -581 101
rect -572 71 -567 101
rect -563 71 -558 101
rect -542 71 -537 101
rect -533 71 -528 101
rect -519 71 -514 101
rect -510 71 -505 101
rect -482 81 -477 111
rect -473 81 -468 111
rect -438 75 -433 105
rect -429 75 -424 105
rect -420 71 -415 101
rect -411 71 -406 101
rect -397 71 -392 101
rect -388 71 -383 101
rect -367 71 -362 101
rect -358 71 -353 101
rect -344 71 -339 101
rect -335 71 -330 101
rect -307 81 -302 111
rect -298 81 -293 111
rect -263 106 -223 111
rect -263 97 -223 102
rect -130 99 -90 104
rect -130 90 -90 95
rect -266 74 -226 79
rect -266 65 -226 70
rect -130 67 -90 72
rect -130 58 -90 63
rect -262 42 -222 47
rect -262 33 -222 38
rect -130 32 -90 37
rect -130 23 -90 28
rect -613 -57 -608 -27
rect -604 -57 -599 -27
rect -595 -61 -590 -31
rect -586 -61 -581 -31
rect -572 -61 -567 -31
rect -563 -61 -558 -31
rect -542 -61 -537 -31
rect -533 -61 -528 -31
rect -519 -61 -514 -31
rect -510 -61 -505 -31
rect -482 -51 -477 -21
rect -473 -51 -468 -21
rect 34 -10 39 30
rect 43 -10 48 30
rect 66 -13 71 27
rect 75 -13 80 27
rect 98 -9 103 31
rect 107 -9 112 31
rect 140 -14 145 46
rect 149 -14 154 46
rect -438 -57 -433 -27
rect -429 -57 -424 -27
rect -420 -61 -415 -31
rect -411 -61 -406 -31
rect -397 -61 -392 -31
rect -388 -61 -383 -31
rect -367 -61 -362 -31
rect -358 -61 -353 -31
rect -344 -61 -339 -31
rect -335 -61 -330 -31
rect -307 -51 -302 -21
rect -298 -51 -293 -21
rect -263 -22 -223 -17
rect 172 -20 177 40
rect 181 -20 186 40
rect 204 -20 209 40
rect 213 -20 218 40
rect 236 7 241 47
rect 245 7 250 47
rect 290 29 295 109
rect 299 29 304 109
rect 464 117 469 157
rect 473 117 478 157
rect 499 116 504 156
rect 508 116 513 156
rect 534 116 539 156
rect 543 116 548 156
rect 569 116 574 156
rect 578 116 583 156
rect 604 116 609 156
rect 613 116 618 156
rect 636 116 641 156
rect 645 116 650 156
rect 773 152 778 182
rect 782 152 787 182
rect 791 148 796 178
rect 800 148 805 178
rect 814 148 819 178
rect 823 148 828 178
rect 844 148 849 178
rect 853 148 858 178
rect 867 148 872 178
rect 876 148 881 178
rect 904 158 909 188
rect 913 158 918 188
rect 322 23 327 103
rect 331 23 336 103
rect 354 23 359 103
rect 363 23 368 103
rect 386 23 391 103
rect 395 23 400 103
rect 418 70 423 110
rect 427 70 432 110
rect -263 -31 -223 -26
rect -130 -29 -90 -24
rect -130 -38 -90 -33
rect -266 -54 -226 -49
rect -266 -63 -226 -58
rect -130 -61 -90 -56
rect -130 -70 -90 -65
rect -262 -86 -222 -81
rect -262 -95 -222 -90
rect -130 -96 -90 -91
rect -130 -105 -90 -100
rect -613 -188 -608 -158
rect -604 -188 -599 -158
rect -595 -192 -590 -162
rect -586 -192 -581 -162
rect -572 -192 -567 -162
rect -563 -192 -558 -162
rect -542 -192 -537 -162
rect -533 -192 -528 -162
rect -519 -192 -514 -162
rect -510 -192 -505 -162
rect -482 -182 -477 -152
rect -473 -182 -468 -152
rect -263 -150 -223 -145
rect -438 -188 -433 -158
rect -429 -188 -424 -158
rect -420 -192 -415 -162
rect -411 -192 -406 -162
rect -397 -192 -392 -162
rect -388 -192 -383 -162
rect -367 -192 -362 -162
rect -358 -192 -353 -162
rect -344 -192 -339 -162
rect -335 -192 -330 -162
rect -307 -182 -302 -152
rect -298 -182 -293 -152
rect -263 -159 -223 -154
rect -130 -157 -90 -152
rect -130 -166 -90 -161
rect 36 -176 41 -116
rect 45 -176 50 -116
rect -266 -182 -226 -177
rect 68 -182 73 -122
rect 77 -182 82 -122
rect 100 -182 105 -122
rect 109 -182 114 -122
rect 132 -155 137 -115
rect 141 -155 146 -115
rect 168 -172 173 -132
rect 177 -172 182 -132
rect 200 -175 205 -135
rect 209 -175 214 -135
rect 232 -171 237 -131
rect 241 -171 246 -131
rect 282 -159 287 -79
rect 291 -159 296 -79
rect 314 -165 319 -85
rect 323 -165 328 -85
rect 346 -165 351 -85
rect 355 -165 360 -85
rect 378 -165 383 -85
rect 387 -165 392 -85
rect 410 -118 415 -78
rect 419 -118 424 -78
rect 451 -85 456 15
rect 460 -85 465 15
rect 668 48 673 88
rect 677 48 682 88
rect 700 48 705 88
rect 709 48 714 88
rect 735 48 740 88
rect 744 48 749 88
rect 773 20 778 50
rect 782 20 787 50
rect 483 -91 488 9
rect 492 -91 497 9
rect 515 -91 520 9
rect 524 -91 529 9
rect 547 -91 552 9
rect 556 -91 561 9
rect 579 -91 584 9
rect 588 -91 593 9
rect 613 -24 618 16
rect 622 -24 627 16
rect 791 16 796 46
rect 800 16 805 46
rect 814 16 819 46
rect 823 16 828 46
rect 844 16 849 46
rect 853 16 858 46
rect 867 16 872 46
rect 876 16 881 46
rect 904 26 909 56
rect 913 26 918 56
rect 668 -97 673 -57
rect 677 -97 682 -57
rect 700 -97 705 -57
rect 709 -97 714 -57
rect 735 -97 740 -57
rect 744 -97 749 -57
rect 773 -111 778 -81
rect 782 -111 787 -81
rect 791 -115 796 -85
rect 800 -115 805 -85
rect 814 -115 819 -85
rect 823 -115 828 -85
rect 844 -115 849 -85
rect 853 -115 858 -85
rect 867 -115 872 -85
rect 876 -115 881 -85
rect 904 -105 909 -75
rect 913 -105 918 -75
rect -266 -191 -226 -186
rect -130 -189 -90 -184
rect -130 -198 -90 -193
rect -262 -214 -222 -209
rect -262 -223 -222 -218
rect -130 -224 -90 -219
rect -130 -233 -90 -228
rect 36 -309 41 -269
rect 45 -309 50 -269
rect 68 -312 73 -272
rect 77 -312 82 -272
rect 100 -308 105 -268
rect 109 -308 114 -268
rect 132 -320 137 -280
rect 141 -320 146 -280
rect 169 -320 174 -280
rect 178 -320 183 -280
rect 201 -319 206 -279
rect 210 -319 215 -279
rect 271 -316 276 -276
rect 280 -316 285 -276
rect 306 -317 311 -277
rect 315 -317 320 -277
rect 341 -317 346 -277
rect 350 -317 355 -277
rect 373 -317 378 -277
rect 382 -317 387 -277
rect 433 -306 438 -266
rect 442 -306 447 -266
rect 645 -244 650 -204
rect 654 -244 659 -204
rect 677 -244 682 -204
rect 686 -244 691 -204
rect 712 -244 717 -204
rect 721 -244 726 -204
rect 773 -243 778 -213
rect 782 -243 787 -213
rect 791 -247 796 -217
rect 800 -247 805 -217
rect 814 -247 819 -217
rect 823 -247 828 -217
rect 844 -247 849 -217
rect 853 -247 858 -217
rect 867 -247 872 -217
rect 876 -247 881 -217
rect 904 -237 909 -207
rect 913 -237 918 -207
rect 468 -307 473 -267
rect 477 -307 482 -267
rect 503 -307 508 -267
rect 512 -307 517 -267
rect 538 -307 543 -267
rect 547 -307 552 -267
rect 570 -307 575 -267
rect 579 -307 584 -267
rect -177 -372 -172 -342
rect -168 -372 -163 -342
rect -159 -376 -154 -346
rect -150 -376 -145 -346
rect -136 -376 -131 -346
rect -127 -376 -122 -346
rect -106 -376 -101 -346
rect -97 -376 -92 -346
rect -83 -376 -78 -346
rect -74 -376 -69 -346
rect -46 -366 -41 -336
rect -37 -366 -32 -336
rect 645 -389 650 -349
rect 654 -389 659 -349
rect 677 -389 682 -349
rect 686 -389 691 -349
rect 712 -389 717 -349
rect 721 -389 726 -349
rect 773 -374 778 -344
rect 782 -374 787 -344
rect 791 -378 796 -348
rect 800 -378 805 -348
rect 814 -378 819 -348
rect 823 -378 828 -348
rect 844 -378 849 -348
rect 853 -378 858 -348
rect 867 -378 872 -348
rect 876 -378 881 -348
rect 904 -368 909 -338
rect 913 -368 918 -338
<< pdcontact >>
rect -613 262 -608 302
rect -604 262 -599 302
rect -578 262 -573 302
rect -569 262 -564 302
rect -546 262 -541 302
rect -537 262 -532 302
rect -514 262 -509 302
rect -505 262 -500 302
rect -482 262 -477 302
rect -473 262 -468 302
rect -438 262 -433 302
rect -429 262 -424 302
rect -403 262 -398 302
rect -394 262 -389 302
rect -371 262 -366 302
rect -362 262 -357 302
rect -339 262 -334 302
rect -330 262 -325 302
rect -307 262 -302 302
rect -298 262 -293 302
rect -195 234 -155 239
rect -195 225 -155 230
rect -63 227 -23 232
rect -63 218 -23 223
rect -195 202 -155 207
rect 26 206 31 246
rect 35 206 40 246
rect 58 206 63 246
rect 67 206 72 246
rect 90 206 95 246
rect 99 206 104 246
rect 137 231 142 271
rect 146 231 151 271
rect 169 231 174 271
rect 178 231 183 271
rect 201 231 206 271
rect 210 231 215 271
rect 233 231 238 271
rect 242 231 247 271
rect -195 193 -155 198
rect -63 195 -23 200
rect -63 186 -23 191
rect -613 131 -608 171
rect -604 131 -599 171
rect -578 131 -573 171
rect -569 131 -564 171
rect -546 131 -541 171
rect -537 131 -532 171
rect -514 131 -509 171
rect -505 131 -500 171
rect -482 131 -477 171
rect -473 131 -468 171
rect -438 131 -433 171
rect -429 131 -424 171
rect -403 131 -398 171
rect -394 131 -389 171
rect -371 131 -366 171
rect -362 131 -357 171
rect -339 131 -334 171
rect -330 131 -325 171
rect -307 131 -302 171
rect -298 131 -293 171
rect -195 170 -155 175
rect -195 161 -155 166
rect -59 160 -19 165
rect -59 151 -19 156
rect 464 198 469 397
rect 473 198 478 397
rect 499 198 504 397
rect 508 198 513 397
rect 534 198 539 397
rect 543 198 548 397
rect 569 198 574 397
rect 578 198 583 397
rect 604 198 609 397
rect 613 198 618 397
rect 290 139 295 179
rect 299 139 304 179
rect 322 139 327 179
rect 331 139 336 179
rect 354 139 359 179
rect 363 139 368 179
rect 386 139 391 179
rect 395 139 400 179
rect 418 139 423 179
rect 427 139 432 179
rect 636 189 641 229
rect 645 189 650 229
rect 773 208 778 248
rect 782 208 787 248
rect 808 208 813 248
rect 817 208 822 248
rect 840 208 845 248
rect 849 208 854 248
rect 872 208 877 248
rect 881 208 886 248
rect 904 208 909 248
rect 913 208 918 248
rect -195 106 -155 111
rect -195 97 -155 102
rect -63 99 -23 104
rect -63 90 -23 95
rect -195 74 -155 79
rect -195 65 -155 70
rect -63 67 -23 72
rect -63 58 -23 63
rect 34 58 39 98
rect 43 58 48 98
rect 66 58 71 98
rect 75 58 80 98
rect 98 58 103 98
rect 107 58 112 98
rect 140 74 145 114
rect 149 74 154 114
rect 172 74 177 114
rect 181 74 186 114
rect 204 74 209 114
rect 213 74 218 114
rect 236 74 241 114
rect 245 74 250 114
rect -195 42 -155 47
rect -613 -1 -608 39
rect -604 -1 -599 39
rect -578 -1 -573 39
rect -569 -1 -564 39
rect -546 -1 -541 39
rect -537 -1 -532 39
rect -514 -1 -509 39
rect -505 -1 -500 39
rect -482 -1 -477 39
rect -473 -1 -468 39
rect -438 -1 -433 39
rect -429 -1 -424 39
rect -403 -1 -398 39
rect -394 -1 -389 39
rect -371 -1 -366 39
rect -362 -1 -357 39
rect -339 -1 -334 39
rect -330 -1 -325 39
rect -307 -1 -302 39
rect -298 -1 -293 39
rect -195 33 -155 38
rect -59 32 -19 37
rect -59 23 -19 28
rect -195 -22 -155 -17
rect 668 115 673 155
rect 677 115 682 155
rect 700 115 705 155
rect 709 115 714 155
rect 735 119 740 159
rect 744 119 749 159
rect 451 51 456 91
rect 460 51 465 91
rect 483 51 488 91
rect 492 51 497 91
rect 515 51 520 91
rect 524 51 529 91
rect 547 51 552 91
rect 556 51 561 91
rect 579 51 584 91
rect 588 51 593 91
rect 613 51 618 91
rect 622 51 627 91
rect -195 -31 -155 -26
rect -63 -29 -23 -24
rect -63 -38 -23 -33
rect -195 -54 -155 -49
rect -195 -63 -155 -58
rect -63 -61 -23 -56
rect -63 -70 -23 -65
rect -195 -86 -155 -81
rect 36 -88 41 -48
rect 45 -88 50 -48
rect 68 -88 73 -48
rect 77 -88 82 -48
rect 100 -88 105 -48
rect 109 -88 114 -48
rect 132 -88 137 -48
rect 141 -88 146 -48
rect 282 -49 287 -9
rect 291 -49 296 -9
rect 314 -49 319 -9
rect 323 -49 328 -9
rect 346 -49 351 -9
rect 355 -49 360 -9
rect 378 -49 383 -9
rect 387 -49 392 -9
rect 410 -49 415 -9
rect 419 -49 424 -9
rect -613 -132 -608 -92
rect -604 -132 -599 -92
rect -578 -132 -573 -92
rect -569 -132 -564 -92
rect -546 -132 -541 -92
rect -537 -132 -532 -92
rect -514 -132 -509 -92
rect -505 -132 -500 -92
rect -482 -132 -477 -92
rect -473 -132 -468 -92
rect -438 -132 -433 -92
rect -429 -132 -424 -92
rect -403 -132 -398 -92
rect -394 -132 -389 -92
rect -371 -132 -366 -92
rect -362 -132 -357 -92
rect -339 -132 -334 -92
rect -330 -132 -325 -92
rect -307 -132 -302 -92
rect -298 -132 -293 -92
rect -195 -95 -155 -90
rect -59 -96 -19 -91
rect -59 -105 -19 -100
rect -195 -150 -155 -145
rect -195 -159 -155 -154
rect -63 -157 -23 -152
rect -63 -166 -23 -161
rect 168 -104 173 -64
rect 177 -104 182 -64
rect 200 -104 205 -64
rect 209 -104 214 -64
rect 232 -104 237 -64
rect 241 -104 246 -64
rect -195 -182 -155 -177
rect 773 76 778 116
rect 782 76 787 116
rect 808 76 813 116
rect 817 76 822 116
rect 840 76 845 116
rect 849 76 854 116
rect 872 76 877 116
rect 881 76 886 116
rect 904 76 909 116
rect 913 76 918 116
rect 668 -30 673 10
rect 677 -30 682 10
rect 700 -30 705 10
rect 709 -30 714 10
rect 735 -26 740 14
rect 744 -26 749 14
rect 773 -55 778 -15
rect 782 -55 787 -15
rect 808 -55 813 -15
rect 817 -55 822 -15
rect 840 -55 845 -15
rect 849 -55 854 -15
rect 872 -55 877 -15
rect 881 -55 886 -15
rect 904 -55 909 -15
rect 913 -55 918 -15
rect -195 -191 -155 -186
rect -63 -189 -23 -184
rect -63 -198 -23 -193
rect -195 -214 -155 -209
rect -195 -223 -155 -218
rect -59 -224 -19 -219
rect -59 -233 -19 -228
rect 36 -241 41 -201
rect 45 -241 50 -201
rect 68 -241 73 -201
rect 77 -241 82 -201
rect 100 -241 105 -201
rect 109 -241 114 -201
rect -177 -316 -172 -276
rect -168 -316 -163 -276
rect -142 -316 -137 -276
rect -133 -316 -128 -276
rect -110 -316 -105 -276
rect -101 -316 -96 -276
rect -78 -316 -73 -276
rect -69 -316 -64 -276
rect -46 -316 -41 -276
rect -37 -316 -32 -276
rect 132 -252 137 -212
rect 141 -252 146 -212
rect 169 -252 174 -212
rect 178 -252 183 -212
rect 201 -252 206 -212
rect 210 -252 215 -212
rect 271 -243 276 -183
rect 280 -243 285 -183
rect 306 -243 311 -183
rect 315 -243 320 -183
rect 341 -243 346 -183
rect 350 -243 355 -183
rect 373 -250 378 -210
rect 382 -250 387 -210
rect 433 -229 438 -149
rect 442 -229 447 -149
rect 468 -229 473 -149
rect 477 -229 482 -149
rect 503 -229 508 -149
rect 512 -229 517 -149
rect 538 -229 543 -149
rect 547 -229 552 -149
rect 645 -177 650 -137
rect 654 -177 659 -137
rect 677 -177 682 -137
rect 686 -177 691 -137
rect 712 -173 717 -133
rect 721 -173 726 -133
rect 570 -236 575 -196
rect 579 -236 584 -196
rect 773 -187 778 -147
rect 782 -187 787 -147
rect 808 -187 813 -147
rect 817 -187 822 -147
rect 840 -187 845 -147
rect 849 -187 854 -147
rect 872 -187 877 -147
rect 881 -187 886 -147
rect 904 -187 909 -147
rect 913 -187 918 -147
rect 645 -322 650 -282
rect 654 -322 659 -282
rect 677 -322 682 -282
rect 686 -322 691 -282
rect 712 -318 717 -278
rect 721 -318 726 -278
rect 773 -318 778 -278
rect 782 -318 787 -278
rect 808 -318 813 -278
rect 817 -318 822 -278
rect 840 -318 845 -278
rect 849 -318 854 -278
rect 872 -318 877 -278
rect 881 -318 886 -278
rect 904 -318 909 -278
rect 913 -318 918 -278
<< polysilicon >>
rect 470 397 472 401
rect 505 397 507 401
rect 540 397 542 401
rect 575 397 577 401
rect 610 397 612 401
rect -607 302 -605 306
rect -572 302 -570 306
rect -540 302 -538 306
rect -508 302 -506 306
rect -476 302 -474 306
rect -432 302 -430 306
rect -397 302 -395 306
rect -365 302 -363 306
rect -333 302 -331 306
rect -301 302 -299 306
rect 143 271 145 275
rect 175 271 177 275
rect 207 271 209 275
rect 239 271 241 275
rect -607 236 -605 262
rect -572 249 -570 262
rect -540 249 -538 262
rect -508 249 -506 262
rect -476 242 -474 262
rect -589 232 -587 240
rect -566 232 -564 240
rect -536 232 -534 240
rect -513 232 -511 240
rect -607 203 -605 206
rect -432 236 -430 262
rect -397 249 -395 262
rect -365 249 -363 262
rect -333 249 -331 262
rect -301 242 -299 262
rect 32 246 34 250
rect 64 246 66 250
rect 96 246 98 250
rect -476 209 -474 212
rect -414 232 -412 240
rect -391 232 -389 240
rect -361 232 -359 240
rect -338 232 -336 240
rect -432 203 -430 206
rect -266 231 -263 233
rect -223 231 -195 233
rect -155 231 -151 233
rect -133 224 -130 226
rect -90 224 -63 226
rect -23 224 -19 226
rect -301 209 -299 212
rect -589 199 -587 202
rect -566 199 -564 202
rect -536 199 -534 202
rect -513 199 -511 202
rect -414 199 -412 202
rect -391 199 -389 202
rect -361 199 -359 202
rect -338 199 -336 202
rect -269 199 -266 201
rect -226 199 -217 201
rect -210 199 -195 201
rect -155 199 -151 201
rect -133 192 -130 194
rect -90 192 -63 194
rect -23 192 -19 194
rect 32 178 34 206
rect 64 191 66 206
rect -607 171 -605 175
rect -572 171 -570 175
rect -540 171 -538 175
rect -508 171 -506 175
rect -476 171 -474 175
rect -432 171 -430 175
rect -397 171 -395 175
rect -365 171 -363 175
rect -333 171 -331 175
rect -301 171 -299 175
rect -265 167 -262 169
rect -222 167 -195 169
rect -155 167 -151 169
rect -133 157 -130 159
rect -90 157 -82 159
rect -75 157 -59 159
rect -19 157 -15 159
rect 64 175 66 184
rect 96 179 98 206
rect 143 203 145 231
rect 175 217 177 231
rect 207 217 209 231
rect 32 135 34 138
rect 175 197 177 205
rect 207 197 209 205
rect 239 204 241 231
rect 143 140 145 143
rect 96 136 98 139
rect 779 248 781 252
rect 814 248 816 252
rect 846 248 848 252
rect 878 248 880 252
rect 910 248 912 252
rect 642 229 644 233
rect 296 179 298 183
rect 328 179 330 183
rect 360 179 362 183
rect 392 179 394 183
rect 424 179 426 183
rect 239 161 241 164
rect 470 157 472 198
rect 505 184 507 198
rect 540 184 542 198
rect 575 184 577 198
rect 610 184 612 198
rect 64 132 66 135
rect 175 133 177 137
rect 207 133 209 137
rect -607 105 -605 131
rect -572 118 -570 131
rect -540 118 -538 131
rect -508 118 -506 131
rect -476 111 -474 131
rect -589 101 -587 109
rect -566 101 -564 109
rect -536 101 -534 109
rect -513 101 -511 109
rect -607 72 -605 75
rect -432 105 -430 131
rect -397 118 -395 131
rect -365 118 -363 131
rect -333 118 -331 131
rect -301 111 -299 131
rect 146 114 148 118
rect 178 114 180 118
rect 210 114 212 118
rect 242 114 244 118
rect -476 78 -474 81
rect -414 101 -412 109
rect -391 101 -389 109
rect -361 101 -359 109
rect -338 101 -336 109
rect -432 72 -430 75
rect -266 103 -263 105
rect -223 103 -195 105
rect -155 103 -151 105
rect 40 98 42 102
rect 72 98 74 102
rect 104 98 106 102
rect -133 96 -130 98
rect -90 96 -63 98
rect -23 96 -19 98
rect -301 78 -299 81
rect -269 71 -266 73
rect -226 71 -217 73
rect -210 71 -195 73
rect -155 71 -151 73
rect -589 68 -587 71
rect -566 68 -564 71
rect -536 68 -534 71
rect -513 68 -511 71
rect -414 68 -412 71
rect -391 68 -389 71
rect -361 68 -359 71
rect -338 68 -336 71
rect -133 64 -130 66
rect -90 64 -63 66
rect -23 64 -19 66
rect 296 109 298 139
rect 328 125 330 139
rect 360 125 362 139
rect 392 125 394 139
rect -607 39 -605 43
rect -572 39 -570 43
rect -540 39 -538 43
rect -508 39 -506 43
rect -476 39 -474 43
rect -432 39 -430 43
rect -397 39 -395 43
rect -365 39 -363 43
rect -333 39 -331 43
rect -301 39 -299 43
rect -265 39 -262 41
rect -222 39 -195 41
rect -155 39 -151 41
rect -133 29 -130 31
rect -90 29 -82 31
rect -75 29 -59 31
rect -19 29 -15 31
rect 40 30 42 58
rect 72 43 74 58
rect -607 -27 -605 -1
rect -572 -14 -570 -1
rect -540 -14 -538 -1
rect -508 -14 -506 -1
rect -476 -21 -474 -1
rect -589 -31 -587 -23
rect -566 -31 -564 -23
rect -536 -31 -534 -23
rect -513 -31 -511 -23
rect -607 -60 -605 -57
rect -432 -27 -430 -1
rect -397 -14 -395 -1
rect -365 -14 -363 -1
rect -333 -14 -331 -1
rect -301 -21 -299 -1
rect 72 27 74 36
rect 104 31 106 58
rect 146 46 148 74
rect 178 60 180 74
rect 210 60 212 74
rect 40 -13 42 -10
rect 104 -12 106 -9
rect 72 -16 74 -13
rect 178 40 180 48
rect 210 40 212 48
rect 242 47 244 74
rect 146 -17 148 -14
rect -476 -54 -474 -51
rect -414 -31 -412 -23
rect -391 -31 -389 -23
rect -361 -31 -359 -23
rect -338 -31 -336 -23
rect -432 -60 -430 -57
rect 328 103 330 111
rect 360 103 362 111
rect 392 103 394 111
rect 424 110 426 139
rect 505 156 507 164
rect 540 156 542 164
rect 575 156 577 164
rect 610 156 612 164
rect 642 156 644 189
rect 779 182 781 208
rect 814 195 816 208
rect 846 195 848 208
rect 878 195 880 208
rect 910 188 912 208
rect 741 159 743 163
rect 470 114 472 117
rect 674 155 676 159
rect 706 155 708 159
rect 505 113 507 116
rect 540 113 542 116
rect 575 113 577 116
rect 610 113 612 116
rect 642 113 644 116
rect 797 178 799 186
rect 820 178 822 186
rect 850 178 852 186
rect 873 178 875 186
rect 779 149 781 152
rect 910 155 912 158
rect 797 145 799 148
rect 820 145 822 148
rect 850 145 852 148
rect 873 145 875 148
rect 296 26 298 29
rect 457 91 459 95
rect 489 91 491 95
rect 521 91 523 95
rect 553 91 555 95
rect 585 91 587 95
rect 619 91 621 95
rect 424 67 426 70
rect 674 88 676 115
rect 706 88 708 115
rect 741 103 743 119
rect 779 116 781 120
rect 814 116 816 120
rect 846 116 848 120
rect 878 116 880 120
rect 910 116 912 120
rect 741 88 743 96
rect 328 19 330 23
rect 360 19 362 23
rect 392 19 394 23
rect 457 15 459 51
rect 489 37 491 51
rect 521 37 523 51
rect 553 37 555 51
rect 585 37 587 51
rect 242 4 244 7
rect 288 -9 290 -5
rect 320 -9 322 -5
rect 352 -9 354 -5
rect 384 -9 386 -5
rect 416 -9 418 -5
rect -266 -25 -263 -23
rect -223 -25 -195 -23
rect -155 -25 -151 -23
rect 178 -24 180 -20
rect 210 -24 212 -20
rect -133 -32 -130 -30
rect -90 -32 -63 -30
rect -23 -32 -19 -30
rect 42 -48 44 -44
rect 74 -48 76 -44
rect 106 -48 108 -44
rect 138 -48 140 -44
rect -301 -54 -299 -51
rect -269 -57 -266 -55
rect -226 -57 -217 -55
rect -210 -57 -195 -55
rect -155 -57 -151 -55
rect -589 -64 -587 -61
rect -566 -64 -564 -61
rect -536 -64 -534 -61
rect -513 -64 -511 -61
rect -414 -64 -412 -61
rect -391 -64 -389 -61
rect -361 -64 -359 -61
rect -338 -64 -336 -61
rect -133 -64 -130 -62
rect -90 -64 -63 -62
rect -23 -64 -19 -62
rect -607 -92 -605 -88
rect -572 -92 -570 -88
rect -540 -92 -538 -88
rect -508 -92 -506 -88
rect -476 -92 -474 -88
rect -432 -92 -430 -88
rect -397 -92 -395 -88
rect -365 -92 -363 -88
rect -333 -92 -331 -88
rect -301 -92 -299 -88
rect -265 -89 -262 -87
rect -222 -89 -195 -87
rect -155 -89 -151 -87
rect 174 -64 176 -60
rect 206 -64 208 -60
rect 238 -64 240 -60
rect -133 -99 -130 -97
rect -90 -99 -82 -97
rect -75 -99 -59 -97
rect -19 -99 -15 -97
rect 42 -116 44 -88
rect 74 -102 76 -88
rect 106 -102 108 -88
rect -607 -158 -605 -132
rect -572 -145 -570 -132
rect -540 -145 -538 -132
rect -508 -145 -506 -132
rect -476 -152 -474 -132
rect -589 -162 -587 -154
rect -566 -162 -564 -154
rect -536 -162 -534 -154
rect -513 -162 -511 -154
rect -607 -191 -605 -188
rect -432 -158 -430 -132
rect -397 -145 -395 -132
rect -365 -145 -363 -132
rect -333 -145 -331 -132
rect -301 -152 -299 -132
rect -476 -185 -474 -182
rect -414 -162 -412 -154
rect -391 -162 -389 -154
rect -361 -162 -359 -154
rect -338 -162 -336 -154
rect -432 -191 -430 -188
rect -266 -153 -263 -151
rect -223 -153 -195 -151
rect -155 -153 -151 -151
rect -133 -160 -130 -158
rect -90 -160 -63 -158
rect -23 -160 -19 -158
rect 74 -122 76 -114
rect 106 -122 108 -114
rect 138 -115 140 -88
rect 288 -79 290 -49
rect 320 -63 322 -49
rect 352 -63 354 -49
rect 384 -63 386 -49
rect -301 -185 -299 -182
rect 42 -179 44 -176
rect 174 -132 176 -104
rect 206 -119 208 -104
rect 138 -158 140 -155
rect 206 -135 208 -126
rect 238 -131 240 -104
rect 174 -175 176 -172
rect 320 -85 322 -77
rect 352 -85 354 -77
rect 384 -85 386 -77
rect 416 -78 418 -49
rect 288 -162 290 -159
rect 489 9 491 17
rect 521 9 523 17
rect 553 9 555 17
rect 585 9 587 17
rect 619 16 621 51
rect 779 50 781 76
rect 814 63 816 76
rect 846 63 848 76
rect 878 63 880 76
rect 910 56 912 76
rect 674 45 676 48
rect 706 45 708 48
rect 741 45 743 48
rect 797 46 799 54
rect 820 46 822 54
rect 850 46 852 54
rect 873 46 875 54
rect 457 -88 459 -85
rect 741 14 743 18
rect 779 17 781 20
rect 910 23 912 26
rect 674 10 676 14
rect 706 10 708 14
rect 619 -27 621 -24
rect 797 13 799 16
rect 820 13 822 16
rect 850 13 852 16
rect 873 13 875 16
rect 779 -15 781 -11
rect 814 -15 816 -11
rect 846 -15 848 -11
rect 878 -15 880 -11
rect 910 -15 912 -11
rect 674 -57 676 -30
rect 706 -57 708 -30
rect 741 -42 743 -26
rect 741 -57 743 -49
rect 489 -95 491 -91
rect 521 -95 523 -91
rect 553 -95 555 -91
rect 585 -95 587 -91
rect 779 -81 781 -55
rect 814 -68 816 -55
rect 846 -68 848 -55
rect 878 -68 880 -55
rect 910 -75 912 -55
rect 674 -100 676 -97
rect 706 -100 708 -97
rect 741 -100 743 -97
rect 797 -85 799 -77
rect 820 -85 822 -77
rect 850 -85 852 -77
rect 873 -85 875 -77
rect 779 -114 781 -111
rect 910 -108 912 -105
rect 797 -118 799 -115
rect 820 -118 822 -115
rect 850 -118 852 -115
rect 873 -118 875 -115
rect 416 -121 418 -118
rect 718 -133 720 -129
rect 651 -137 653 -133
rect 683 -137 685 -133
rect 439 -149 441 -145
rect 474 -149 476 -145
rect 509 -149 511 -145
rect 544 -149 546 -145
rect 320 -169 322 -165
rect 352 -169 354 -165
rect 384 -169 386 -165
rect 238 -174 240 -171
rect 206 -178 208 -175
rect -269 -185 -266 -183
rect -226 -185 -217 -183
rect -210 -185 -195 -183
rect -155 -185 -151 -183
rect 74 -186 76 -182
rect 106 -186 108 -182
rect 277 -183 279 -179
rect 312 -183 314 -179
rect 347 -183 349 -179
rect -133 -192 -130 -190
rect -90 -192 -63 -190
rect -23 -192 -19 -190
rect -589 -195 -587 -192
rect -566 -195 -564 -192
rect -536 -195 -534 -192
rect -513 -195 -511 -192
rect -414 -195 -412 -192
rect -391 -195 -389 -192
rect -361 -195 -359 -192
rect -338 -195 -336 -192
rect 42 -201 44 -197
rect 74 -201 76 -197
rect 106 -201 108 -197
rect -265 -217 -262 -215
rect -222 -217 -195 -215
rect -155 -217 -151 -215
rect -133 -227 -130 -225
rect -90 -227 -82 -225
rect -75 -227 -59 -225
rect -19 -227 -15 -225
rect 138 -212 140 -208
rect 175 -212 177 -208
rect 207 -212 209 -208
rect 42 -269 44 -241
rect 74 -256 76 -241
rect -171 -276 -169 -272
rect -136 -276 -134 -272
rect -104 -276 -102 -272
rect -72 -276 -70 -272
rect -40 -276 -38 -272
rect 74 -272 76 -263
rect 106 -268 108 -241
rect 379 -210 381 -206
rect 42 -312 44 -309
rect 138 -280 140 -252
rect 175 -280 177 -252
rect 207 -279 209 -252
rect 277 -276 279 -243
rect 312 -257 314 -243
rect 347 -257 349 -243
rect 779 -147 781 -143
rect 814 -147 816 -143
rect 846 -147 848 -143
rect 878 -147 880 -143
rect 910 -147 912 -143
rect 576 -196 578 -192
rect 106 -311 108 -308
rect 74 -315 76 -312
rect -171 -342 -169 -316
rect -136 -329 -134 -316
rect -104 -329 -102 -316
rect -72 -329 -70 -316
rect -40 -336 -38 -316
rect 312 -277 314 -269
rect 347 -277 349 -269
rect 379 -277 381 -250
rect 439 -266 441 -229
rect 474 -243 476 -229
rect 509 -243 511 -229
rect 544 -243 546 -229
rect 651 -204 653 -177
rect 683 -204 685 -177
rect 718 -189 720 -173
rect 718 -204 720 -196
rect 277 -319 279 -316
rect 474 -267 476 -259
rect 509 -267 511 -259
rect 544 -267 546 -259
rect 576 -267 578 -236
rect 779 -213 781 -187
rect 814 -200 816 -187
rect 846 -200 848 -187
rect 878 -200 880 -187
rect 910 -207 912 -187
rect 797 -217 799 -209
rect 820 -217 822 -209
rect 850 -217 852 -209
rect 873 -217 875 -209
rect 651 -247 653 -244
rect 683 -247 685 -244
rect 718 -247 720 -244
rect 779 -246 781 -243
rect 910 -240 912 -237
rect 797 -250 799 -247
rect 820 -250 822 -247
rect 850 -250 852 -247
rect 873 -250 875 -247
rect 439 -309 441 -306
rect 718 -278 720 -274
rect 779 -278 781 -274
rect 814 -278 816 -274
rect 846 -278 848 -274
rect 878 -278 880 -274
rect 910 -278 912 -274
rect 651 -282 653 -278
rect 683 -282 685 -278
rect 474 -310 476 -307
rect 509 -310 511 -307
rect 544 -310 546 -307
rect 576 -310 578 -307
rect 138 -323 140 -320
rect 175 -323 177 -320
rect 207 -322 209 -319
rect 312 -320 314 -317
rect 347 -320 349 -317
rect 379 -320 381 -317
rect -153 -346 -151 -338
rect -130 -346 -128 -338
rect -100 -346 -98 -338
rect -77 -346 -75 -338
rect -171 -375 -169 -372
rect 651 -349 653 -322
rect 683 -349 685 -322
rect 718 -334 720 -318
rect 718 -349 720 -341
rect 779 -344 781 -318
rect 814 -331 816 -318
rect 846 -331 848 -318
rect 878 -331 880 -318
rect 910 -338 912 -318
rect -40 -369 -38 -366
rect -153 -379 -151 -376
rect -130 -379 -128 -376
rect -100 -379 -98 -376
rect -77 -379 -75 -376
rect 797 -348 799 -340
rect 820 -348 822 -340
rect 850 -348 852 -340
rect 873 -348 875 -340
rect 779 -377 781 -374
rect 910 -371 912 -368
rect 797 -381 799 -378
rect 820 -381 822 -378
rect 850 -381 852 -378
rect 873 -381 875 -378
rect 651 -392 653 -389
rect 683 -392 685 -389
rect 718 -392 720 -389
<< polycontact >>
rect -612 239 -607 243
rect -577 249 -572 254
rect -545 249 -540 254
rect -513 249 -508 254
rect -481 245 -476 250
rect -594 235 -589 240
rect -571 235 -566 240
rect -541 235 -536 240
rect -518 235 -513 240
rect -437 239 -432 243
rect -402 249 -397 254
rect -370 249 -365 254
rect -338 249 -333 254
rect -306 245 -301 250
rect -419 235 -414 240
rect -396 235 -391 240
rect -366 235 -361 240
rect -343 235 -338 240
rect -209 233 -204 238
rect -77 226 -72 231
rect -223 201 -218 206
rect -209 201 -204 206
rect 138 217 143 222
rect -86 194 -81 199
rect 27 192 32 197
rect 59 192 64 197
rect 91 187 96 192
rect 59 178 64 183
rect -214 169 -209 174
rect -87 159 -83 163
rect -72 159 -67 164
rect 170 217 175 222
rect 202 217 207 222
rect 234 210 239 215
rect 170 200 175 205
rect 202 200 207 205
rect 465 181 470 186
rect 500 184 505 189
rect 535 184 540 189
rect 570 184 575 189
rect 605 184 610 189
rect 637 173 642 178
rect 500 159 505 164
rect -612 108 -607 112
rect -577 118 -572 123
rect -545 118 -540 123
rect -513 118 -508 123
rect -481 114 -476 119
rect -594 104 -589 109
rect -571 104 -566 109
rect -541 104 -536 109
rect -518 104 -513 109
rect -437 108 -432 112
rect -402 118 -397 123
rect -370 118 -365 123
rect -338 118 -333 123
rect -306 114 -301 119
rect 291 125 296 130
rect -419 104 -414 109
rect -396 104 -391 109
rect -366 104 -361 109
rect -343 104 -338 109
rect -209 105 -204 110
rect -77 98 -72 103
rect -223 73 -218 78
rect -209 73 -204 78
rect -86 66 -81 71
rect 323 125 328 130
rect 355 125 360 130
rect 387 125 392 130
rect 419 118 424 123
rect 141 60 146 65
rect -214 41 -209 46
rect 35 44 40 49
rect -87 31 -83 35
rect -72 31 -67 36
rect 67 44 72 49
rect 99 39 104 44
rect 67 30 72 35
rect -612 -24 -607 -20
rect -577 -14 -572 -9
rect -545 -14 -540 -9
rect -513 -14 -508 -9
rect -481 -18 -476 -13
rect -594 -28 -589 -23
rect -571 -28 -566 -23
rect -541 -28 -536 -23
rect -518 -28 -513 -23
rect -437 -24 -432 -20
rect -402 -14 -397 -9
rect -370 -14 -365 -9
rect -338 -14 -333 -9
rect -306 -18 -301 -13
rect 173 60 178 65
rect 205 60 210 65
rect 237 53 242 58
rect 173 43 178 48
rect 205 43 210 48
rect -419 -28 -414 -23
rect -396 -28 -391 -23
rect -366 -28 -361 -23
rect -343 -28 -338 -23
rect -209 -23 -204 -18
rect 323 106 328 111
rect 355 106 360 111
rect 387 106 392 111
rect 535 159 540 164
rect 570 159 575 164
rect 605 159 610 164
rect 774 185 779 189
rect 809 195 814 200
rect 841 195 846 200
rect 873 195 878 200
rect 905 191 910 196
rect 792 181 797 186
rect 815 181 820 186
rect 845 181 850 186
rect 868 181 873 186
rect 669 101 674 106
rect 701 92 706 97
rect 736 106 741 111
rect 737 91 741 95
rect 452 37 457 42
rect 484 37 489 42
rect 516 37 521 42
rect 548 37 553 42
rect 580 37 585 42
rect 614 30 619 35
rect -77 -30 -72 -25
rect -223 -55 -218 -50
rect -209 -55 -204 -50
rect -86 -62 -81 -57
rect -214 -87 -209 -82
rect 283 -63 288 -58
rect -87 -97 -83 -93
rect -72 -97 -67 -92
rect 37 -102 42 -97
rect 69 -102 74 -97
rect 101 -102 106 -97
rect 133 -109 138 -104
rect -612 -155 -607 -151
rect -577 -145 -572 -140
rect -545 -145 -540 -140
rect -513 -145 -508 -140
rect -481 -149 -476 -144
rect -594 -159 -589 -154
rect -571 -159 -566 -154
rect -541 -159 -536 -154
rect -518 -159 -513 -154
rect -437 -155 -432 -151
rect -402 -145 -397 -140
rect -370 -145 -365 -140
rect -338 -145 -333 -140
rect -306 -149 -301 -144
rect -209 -151 -204 -146
rect -419 -159 -414 -154
rect -396 -159 -391 -154
rect -366 -159 -361 -154
rect -343 -159 -338 -154
rect -77 -158 -72 -153
rect 69 -119 74 -114
rect 101 -119 106 -114
rect 315 -63 320 -58
rect 347 -63 352 -58
rect 379 -63 384 -58
rect 411 -70 416 -65
rect -223 -183 -218 -178
rect -209 -183 -204 -178
rect 169 -118 174 -113
rect 201 -118 206 -113
rect 233 -123 238 -118
rect 201 -132 206 -127
rect 315 -82 320 -77
rect 347 -82 352 -77
rect 379 -82 384 -77
rect 484 12 489 17
rect 516 12 521 17
rect 548 12 553 17
rect 580 12 585 17
rect 774 53 779 57
rect 809 63 814 68
rect 841 63 846 68
rect 873 63 878 68
rect 905 59 910 64
rect 792 49 797 54
rect 815 49 820 54
rect 845 49 850 54
rect 868 49 873 54
rect 669 -44 674 -39
rect 701 -53 706 -48
rect 736 -39 741 -34
rect 737 -54 741 -50
rect 774 -78 779 -74
rect 809 -68 814 -63
rect 841 -68 846 -63
rect 873 -68 878 -63
rect 905 -72 910 -67
rect 792 -82 797 -77
rect 815 -82 820 -77
rect 845 -82 850 -77
rect 868 -82 873 -77
rect -86 -190 -81 -185
rect -214 -215 -209 -210
rect -87 -225 -83 -221
rect -72 -225 -67 -220
rect 37 -255 42 -250
rect 69 -255 74 -250
rect 101 -260 106 -255
rect 69 -269 74 -264
rect 133 -266 138 -261
rect 170 -266 175 -261
rect 202 -271 207 -266
rect 272 -260 277 -255
rect 307 -257 312 -252
rect 342 -257 347 -252
rect 646 -191 651 -186
rect 434 -246 439 -241
rect 307 -274 312 -269
rect -176 -339 -171 -335
rect -141 -329 -136 -324
rect -109 -329 -104 -324
rect -77 -329 -72 -324
rect -45 -333 -40 -328
rect 342 -274 347 -269
rect 374 -271 379 -266
rect 469 -243 474 -238
rect 504 -243 509 -238
rect 539 -243 544 -238
rect 678 -200 683 -195
rect 713 -186 718 -181
rect 714 -201 718 -197
rect 571 -252 576 -247
rect 469 -264 474 -259
rect 504 -264 509 -259
rect 539 -264 544 -259
rect 774 -210 779 -206
rect 809 -200 814 -195
rect 841 -200 846 -195
rect 873 -200 878 -195
rect 905 -204 910 -199
rect 792 -214 797 -209
rect 815 -214 820 -209
rect 845 -214 850 -209
rect 868 -214 873 -209
rect 646 -336 651 -331
rect -158 -343 -153 -338
rect -135 -343 -130 -338
rect -105 -343 -100 -338
rect -82 -343 -77 -338
rect 678 -345 683 -340
rect 713 -331 718 -326
rect 774 -341 779 -337
rect 714 -346 718 -342
rect 809 -331 814 -326
rect 841 -331 846 -326
rect 873 -331 878 -326
rect 905 -335 910 -330
rect 792 -345 797 -340
rect 815 -345 820 -340
rect 845 -345 850 -340
rect 868 -345 873 -340
<< metal1 >>
rect 458 403 484 406
rect 487 403 519 406
rect 522 403 554 406
rect 557 403 589 406
rect 592 403 624 406
rect 464 397 469 403
rect -613 314 -564 317
rect -438 314 -389 317
rect -613 302 -608 314
rect -567 311 -477 314
rect -590 308 -573 311
rect -604 256 -599 262
rect -590 256 -587 308
rect -578 302 -573 308
rect -546 302 -541 311
rect -514 302 -509 311
rect -482 302 -477 311
rect -438 302 -433 314
rect -392 311 -302 314
rect -415 308 -398 311
rect -604 253 -587 256
rect -579 249 -577 254
rect -604 246 -583 249
rect -569 246 -564 262
rect -537 254 -532 262
rect -547 249 -545 254
rect -537 249 -513 254
rect -505 250 -500 262
rect -473 253 -468 262
rect -429 256 -424 262
rect -415 256 -412 308
rect -403 302 -398 308
rect -371 302 -366 311
rect -339 302 -334 311
rect -307 302 -302 311
rect -429 253 -412 256
rect -473 250 -454 253
rect -537 246 -532 249
rect -619 239 -612 243
rect -604 236 -599 246
rect -586 243 -564 246
rect -558 243 -532 246
rect -505 245 -481 250
rect -594 240 -589 242
rect -571 240 -566 243
rect -586 233 -575 236
rect -558 238 -554 243
rect -563 235 -554 238
rect -541 240 -536 243
rect -518 240 -513 242
rect -586 232 -581 233
rect -613 202 -608 206
rect -578 202 -575 233
rect -563 232 -558 235
rect -533 233 -522 236
rect -505 238 -500 245
rect -473 242 -468 250
rect -404 249 -402 254
rect -429 246 -408 249
rect -394 246 -389 262
rect -362 254 -357 262
rect -372 249 -370 254
rect -362 249 -338 254
rect -330 250 -325 262
rect -298 251 -293 262
rect 118 283 265 286
rect 20 252 110 258
rect -362 246 -357 249
rect -510 235 -500 238
rect -533 232 -528 233
rect -525 202 -522 233
rect -510 232 -505 235
rect -443 239 -437 243
rect -429 236 -424 246
rect -411 243 -389 246
rect -383 243 -357 246
rect -330 245 -306 250
rect -298 246 -287 251
rect 26 246 31 252
rect 58 246 63 252
rect 90 246 95 252
rect -613 199 -590 202
rect -578 199 -567 202
rect -594 196 -590 199
rect -542 196 -537 202
rect -525 199 -514 202
rect -482 196 -477 212
rect -419 240 -414 242
rect -396 240 -391 243
rect -411 233 -400 236
rect -383 238 -379 243
rect -388 235 -379 238
rect -366 240 -361 243
rect -343 240 -338 242
rect -411 232 -406 233
rect -438 202 -433 206
rect -403 202 -400 233
rect -388 232 -383 235
rect -358 233 -347 236
rect -330 238 -325 245
rect -298 242 -293 246
rect -335 235 -325 238
rect -358 232 -353 233
rect -350 202 -347 233
rect -335 232 -330 235
rect -277 234 -263 239
rect -209 238 -204 244
rect -438 199 -415 202
rect -403 199 -392 202
rect -594 193 -477 196
rect -419 196 -415 199
rect -367 196 -362 202
rect -350 199 -339 202
rect -307 196 -302 212
rect -419 193 -302 196
rect -613 183 -564 186
rect -438 183 -389 186
rect -613 171 -608 183
rect -567 180 -477 183
rect -590 177 -573 180
rect -604 125 -599 131
rect -590 125 -587 177
rect -578 171 -573 177
rect -546 171 -541 180
rect -514 171 -509 180
rect -482 171 -477 180
rect -438 171 -433 183
rect -392 180 -302 183
rect -415 177 -398 180
rect -604 122 -587 125
rect -579 118 -577 123
rect -604 115 -583 118
rect -569 115 -564 131
rect -537 123 -532 131
rect -547 118 -545 123
rect -537 118 -513 123
rect -505 119 -500 131
rect -473 122 -468 131
rect -429 125 -424 131
rect -415 125 -412 177
rect -403 171 -398 177
rect -371 171 -366 180
rect -339 171 -334 180
rect -307 171 -302 180
rect -277 175 -273 234
rect -155 234 -143 239
rect -223 222 -219 230
rect -270 218 -219 222
rect -209 225 -195 230
rect -209 219 -204 225
rect -270 202 -266 218
rect -215 214 -204 219
rect -223 206 -218 209
rect -215 198 -212 214
rect -209 206 -204 209
rect -149 207 -143 234
rect -140 227 -130 232
rect -77 231 -72 237
rect -17 232 -11 238
rect -140 218 -136 227
rect -23 227 -11 232
rect -90 218 -63 223
rect -77 212 -72 218
rect -17 212 -11 227
rect -155 202 -143 207
rect -226 193 -195 198
rect -277 170 -262 175
rect -214 174 -209 193
rect -149 175 -143 202
rect -140 207 -72 212
rect -140 200 -137 207
rect -140 195 -130 200
rect -86 199 -81 202
rect -140 179 -137 195
rect -23 195 -12 200
rect 35 197 40 206
rect 23 192 27 197
rect 35 192 51 197
rect 56 192 59 197
rect 67 192 72 206
rect 99 192 104 206
rect 118 192 121 283
rect 131 277 253 280
rect 137 271 142 277
rect 169 271 174 277
rect 201 271 206 277
rect 233 271 238 277
rect 124 217 138 222
rect 146 213 151 231
rect 167 217 170 222
rect 178 213 183 231
rect 199 217 202 222
rect 210 213 215 231
rect 242 217 247 231
rect 227 213 234 215
rect 146 210 234 213
rect 242 212 250 217
rect 146 203 160 207
rect -90 186 -63 191
rect 46 189 51 192
rect 67 189 91 192
rect 46 187 91 189
rect 99 187 121 192
rect 46 186 72 187
rect -140 175 -83 179
rect -155 170 -143 175
rect -222 161 -195 166
rect -214 139 -209 161
rect -135 160 -130 165
rect -87 163 -83 175
rect -80 156 -77 186
rect 35 178 47 182
rect 56 178 59 183
rect -72 164 -67 167
rect -19 160 -8 165
rect -90 151 -59 156
rect -77 145 -72 151
rect -429 122 -412 125
rect -473 119 -454 122
rect -537 115 -532 118
rect -619 108 -612 112
rect -604 105 -599 115
rect -586 112 -564 115
rect -558 112 -532 115
rect -505 114 -481 119
rect -594 109 -589 111
rect -571 109 -566 112
rect -586 102 -575 105
rect -558 107 -554 112
rect -563 104 -554 107
rect -541 109 -536 112
rect -518 109 -513 111
rect -586 101 -581 102
rect -613 71 -608 75
rect -578 71 -575 102
rect -563 101 -558 104
rect -533 102 -522 105
rect -505 107 -500 114
rect -473 111 -468 119
rect -404 118 -402 123
rect -429 115 -408 118
rect -394 115 -389 131
rect -362 123 -357 131
rect -372 118 -370 123
rect -362 118 -338 123
rect -330 119 -325 131
rect -298 122 -293 131
rect 26 128 31 138
rect 43 135 47 178
rect 67 175 72 186
rect 99 179 104 187
rect 137 139 142 143
rect 43 131 63 135
rect 90 128 95 139
rect 137 133 151 139
rect 156 137 160 203
rect 167 200 170 205
rect 178 197 194 201
rect 199 200 202 205
rect 210 197 215 210
rect 242 204 247 212
rect 190 137 194 197
rect 262 199 265 283
rect 439 209 442 210
rect 439 206 456 209
rect 439 205 442 206
rect 262 196 449 199
rect 284 185 438 188
rect 290 179 295 185
rect 322 179 327 185
rect 354 179 359 185
rect 386 179 391 185
rect 418 179 423 185
rect 233 157 238 164
rect 233 153 247 157
rect 446 161 449 196
rect 453 186 456 206
rect 473 188 478 198
rect 487 188 490 403
rect 499 397 504 403
rect 453 181 465 186
rect 473 185 490 188
rect 497 184 500 189
rect 508 188 513 198
rect 522 188 525 403
rect 534 397 539 403
rect 508 185 525 188
rect 532 184 535 189
rect 543 188 548 198
rect 557 188 560 403
rect 569 397 574 403
rect 543 185 560 188
rect 564 184 570 189
rect 578 188 583 198
rect 592 188 595 403
rect 604 397 609 403
rect 773 260 822 263
rect 773 248 778 260
rect 819 257 909 260
rect 796 254 813 257
rect 630 235 656 238
rect 578 185 595 188
rect 602 184 605 189
rect 613 179 618 198
rect 636 229 641 235
rect 782 202 787 208
rect 796 202 799 254
rect 808 248 813 254
rect 840 248 845 257
rect 872 248 877 257
rect 904 248 909 257
rect 782 199 799 202
rect 807 195 809 200
rect 782 192 803 195
rect 817 192 822 208
rect 849 200 854 208
rect 839 195 841 200
rect 849 195 873 200
rect 881 196 886 208
rect 913 199 918 208
rect 913 196 924 199
rect 849 192 854 195
rect 473 178 618 179
rect 645 181 650 189
rect 673 185 774 189
rect 673 181 678 185
rect 782 182 787 192
rect 800 189 822 192
rect 828 189 854 192
rect 881 191 905 196
rect 473 176 637 178
rect 473 157 478 176
rect 497 159 500 164
rect 156 133 174 137
rect 190 133 206 137
rect 26 124 95 128
rect 278 125 291 130
rect -362 115 -357 118
rect -510 104 -500 107
rect -533 101 -528 102
rect -525 71 -522 102
rect -510 101 -505 104
rect -443 108 -437 112
rect -429 105 -424 115
rect -411 112 -389 115
rect -383 112 -357 115
rect -330 114 -306 119
rect -298 117 -287 122
rect 134 120 256 123
rect 299 122 304 139
rect 320 125 323 130
rect 331 122 336 139
rect 352 125 355 130
rect 363 122 368 139
rect 384 125 387 130
rect 395 123 400 139
rect 427 125 432 139
rect 449 125 454 128
rect 395 122 419 123
rect -613 68 -590 71
rect -578 68 -567 71
rect -594 65 -590 68
rect -542 65 -537 71
rect -525 68 -514 71
rect -482 65 -477 81
rect -419 109 -414 111
rect -396 109 -391 112
rect -411 102 -400 105
rect -383 107 -379 112
rect -388 104 -379 107
rect -366 109 -361 112
rect -343 109 -338 111
rect -411 101 -406 102
rect -438 71 -433 75
rect -403 71 -400 102
rect -388 101 -383 104
rect -358 102 -347 105
rect -330 107 -325 114
rect -298 111 -293 117
rect -335 104 -325 107
rect -358 101 -353 102
rect -350 71 -347 102
rect -335 101 -330 104
rect -277 106 -263 111
rect -209 110 -204 116
rect 140 114 145 120
rect 172 114 177 120
rect 204 114 209 120
rect 236 114 241 120
rect 299 119 419 122
rect 395 118 419 119
rect 427 120 454 125
rect -438 68 -415 71
rect -403 68 -392 71
rect -594 62 -477 65
rect -419 65 -415 68
rect -367 65 -362 71
rect -350 68 -339 71
rect -307 65 -302 81
rect -419 62 -302 65
rect -613 51 -564 54
rect -438 51 -389 54
rect -613 39 -608 51
rect -567 48 -477 51
rect -590 45 -573 48
rect -604 -7 -599 -1
rect -590 -7 -587 45
rect -578 39 -573 45
rect -546 39 -541 48
rect -514 39 -509 48
rect -482 39 -477 48
rect -438 39 -433 51
rect -392 48 -302 51
rect -415 45 -398 48
rect -604 -10 -587 -7
rect -579 -14 -577 -9
rect -604 -17 -583 -14
rect -569 -17 -564 -1
rect -537 -9 -532 -1
rect -547 -14 -545 -9
rect -537 -14 -513 -9
rect -505 -13 -500 -1
rect -473 -10 -468 -1
rect -429 -7 -424 -1
rect -415 -7 -412 45
rect -403 39 -398 45
rect -371 39 -366 48
rect -339 39 -334 48
rect -307 39 -302 48
rect -277 47 -273 106
rect -155 110 -149 111
rect -155 106 -143 110
rect -223 94 -219 102
rect -270 90 -219 94
rect -209 97 -195 102
rect -209 91 -204 97
rect -270 74 -266 90
rect -215 86 -204 91
rect -223 78 -218 81
rect -215 70 -212 86
rect -209 78 -204 81
rect -149 79 -143 106
rect -140 99 -130 104
rect -77 103 -72 109
rect -17 104 -11 110
rect 28 104 118 110
rect -140 90 -136 99
rect -23 99 -11 104
rect -90 90 -63 95
rect -77 84 -72 90
rect -17 84 -11 99
rect 34 98 39 104
rect 66 98 71 104
rect 98 98 103 104
rect -155 74 -143 79
rect -226 65 -195 70
rect -277 42 -262 47
rect -214 46 -209 65
rect -149 47 -143 74
rect -140 79 -72 84
rect -140 72 -137 79
rect -140 67 -130 72
rect -86 71 -81 74
rect -140 51 -137 67
rect -23 67 -12 72
rect -90 58 -63 63
rect 299 109 313 112
rect 119 60 141 65
rect -140 47 -83 51
rect -155 42 -143 47
rect -149 41 -143 42
rect -222 33 -195 38
rect -214 11 -209 33
rect -135 32 -130 37
rect -87 35 -83 47
rect -80 28 -77 58
rect 43 49 48 58
rect 17 44 35 49
rect 43 44 59 49
rect 64 44 67 49
rect 75 44 80 58
rect 107 44 112 58
rect 149 56 154 74
rect 170 60 173 65
rect 181 56 186 74
rect 202 60 205 65
rect 213 56 218 74
rect 245 60 250 74
rect 230 56 237 58
rect 149 53 237 56
rect 245 55 267 60
rect 149 46 163 50
rect 54 41 59 44
rect 75 41 99 44
rect 54 39 99 41
rect 107 39 119 44
rect -72 36 -67 39
rect 54 38 80 39
rect -19 32 -8 37
rect 43 30 55 34
rect 64 30 67 35
rect -90 23 -59 28
rect -77 17 -72 23
rect -429 -10 -412 -7
rect -473 -13 -454 -10
rect -537 -17 -532 -14
rect -619 -24 -612 -20
rect -604 -27 -599 -17
rect -586 -20 -564 -17
rect -558 -20 -532 -17
rect -505 -18 -481 -13
rect -594 -23 -589 -21
rect -571 -23 -566 -20
rect -586 -30 -575 -27
rect -558 -25 -554 -20
rect -563 -28 -554 -25
rect -541 -23 -536 -20
rect -518 -23 -513 -21
rect -586 -31 -581 -30
rect -613 -61 -608 -57
rect -578 -61 -575 -30
rect -563 -31 -558 -28
rect -533 -30 -522 -27
rect -505 -25 -500 -18
rect -473 -21 -468 -13
rect -404 -14 -402 -9
rect -429 -17 -408 -14
rect -394 -17 -389 -1
rect -362 -9 -357 -1
rect -372 -14 -370 -9
rect -362 -14 -338 -9
rect -330 -13 -325 -1
rect -298 -10 -293 -1
rect -362 -17 -357 -14
rect -510 -28 -500 -25
rect -533 -31 -528 -30
rect -525 -61 -522 -30
rect -510 -31 -505 -28
rect -443 -24 -437 -20
rect -429 -27 -424 -17
rect -411 -20 -389 -17
rect -383 -20 -357 -17
rect -330 -18 -306 -13
rect -298 -15 -287 -10
rect -613 -64 -590 -61
rect -578 -64 -567 -61
rect -594 -67 -590 -64
rect -542 -67 -537 -61
rect -525 -64 -514 -61
rect -482 -67 -477 -51
rect -419 -23 -414 -21
rect -396 -23 -391 -20
rect -411 -30 -400 -27
rect -383 -25 -379 -20
rect -388 -28 -379 -25
rect -366 -23 -361 -20
rect -343 -23 -338 -21
rect -411 -31 -406 -30
rect -438 -61 -433 -57
rect -403 -61 -400 -30
rect -388 -31 -383 -28
rect -358 -30 -347 -27
rect -330 -25 -325 -18
rect -298 -21 -293 -15
rect -335 -28 -325 -25
rect -358 -31 -353 -30
rect -350 -61 -347 -30
rect -335 -31 -330 -28
rect -277 -22 -263 -17
rect -209 -18 -204 -12
rect -149 -17 -143 -11
rect -438 -64 -415 -61
rect -403 -64 -392 -61
rect -594 -70 -477 -67
rect -419 -67 -415 -64
rect -367 -67 -362 -61
rect -350 -64 -339 -61
rect -307 -67 -302 -51
rect -419 -70 -302 -67
rect -613 -80 -564 -77
rect -438 -80 -389 -77
rect -613 -92 -608 -80
rect -567 -83 -477 -80
rect -590 -86 -573 -83
rect -604 -138 -599 -132
rect -590 -138 -587 -86
rect -578 -92 -573 -86
rect -546 -92 -541 -83
rect -514 -92 -509 -83
rect -482 -92 -477 -83
rect -438 -92 -433 -80
rect -392 -83 -302 -80
rect -415 -86 -398 -83
rect -604 -141 -587 -138
rect -579 -145 -577 -140
rect -604 -148 -583 -145
rect -569 -148 -564 -132
rect -537 -140 -532 -132
rect -547 -145 -545 -140
rect -537 -145 -513 -140
rect -505 -144 -500 -132
rect -473 -141 -468 -132
rect -429 -138 -424 -132
rect -415 -138 -412 -86
rect -403 -92 -398 -86
rect -371 -92 -366 -83
rect -339 -92 -334 -83
rect -307 -92 -302 -83
rect -277 -81 -273 -22
rect -155 -22 -143 -17
rect -223 -34 -219 -26
rect -270 -38 -219 -34
rect -209 -31 -195 -26
rect -209 -37 -204 -31
rect -270 -54 -266 -38
rect -215 -42 -204 -37
rect -223 -50 -218 -47
rect -215 -58 -212 -42
rect -209 -50 -204 -47
rect -149 -49 -143 -22
rect -140 -29 -130 -24
rect -77 -25 -72 -19
rect -17 -24 -11 -18
rect 34 -20 39 -10
rect 51 -13 55 30
rect 75 27 80 38
rect 107 31 112 39
rect 51 -17 71 -13
rect 98 -20 103 -9
rect 34 -24 103 -20
rect -140 -38 -136 -29
rect -23 -29 -11 -24
rect -90 -38 -63 -33
rect -77 -44 -72 -38
rect -17 -44 -11 -29
rect 116 -27 119 39
rect 140 -18 145 -14
rect 140 -24 154 -18
rect 159 -20 163 46
rect 170 43 173 48
rect 181 40 197 44
rect 202 43 205 48
rect 213 40 218 53
rect 245 47 250 55
rect 193 -20 197 40
rect 262 28 267 55
rect 290 25 295 29
rect 290 19 304 25
rect 309 23 313 109
rect 320 106 323 111
rect 331 103 347 107
rect 352 106 355 111
rect 363 103 379 107
rect 384 106 387 111
rect 395 103 400 118
rect 427 110 432 120
rect 343 23 347 103
rect 375 23 379 103
rect 508 156 513 176
rect 532 159 535 164
rect 543 156 548 176
rect 578 175 637 176
rect 564 159 570 164
rect 578 156 583 175
rect 613 173 637 175
rect 645 176 678 181
rect 602 159 605 164
rect 613 156 618 173
rect 645 156 650 176
rect 662 161 688 167
rect 464 112 469 117
rect 668 155 673 161
rect 700 155 705 166
rect 735 159 740 170
rect 499 112 504 116
rect 534 112 539 116
rect 569 112 574 116
rect 604 112 609 116
rect 636 112 641 116
rect 792 186 797 188
rect 815 186 820 189
rect 800 179 811 182
rect 828 184 832 189
rect 823 181 832 184
rect 845 186 850 189
rect 868 186 873 188
rect 800 178 805 179
rect 773 148 778 152
rect 808 148 811 179
rect 823 178 828 181
rect 853 179 864 182
rect 881 184 886 191
rect 913 188 918 196
rect 876 181 886 184
rect 853 178 858 179
rect 861 148 864 179
rect 876 178 881 181
rect 773 145 796 148
rect 808 145 819 148
rect 792 142 796 145
rect 844 142 849 148
rect 861 145 872 148
rect 904 142 909 158
rect 792 139 909 142
rect 464 109 641 112
rect 455 106 461 109
rect 677 106 682 115
rect 455 103 641 106
rect 445 97 633 100
rect 451 91 456 97
rect 483 91 488 97
rect 515 91 520 97
rect 547 91 552 97
rect 579 91 584 97
rect 613 91 618 97
rect 418 63 423 70
rect 418 59 432 63
rect 439 42 444 45
rect 439 37 452 42
rect 460 34 465 51
rect 481 37 484 42
rect 492 34 497 51
rect 513 37 516 42
rect 524 34 529 51
rect 545 37 548 42
rect 556 34 561 51
rect 577 37 580 42
rect 588 35 593 51
rect 622 37 627 51
rect 638 37 641 103
rect 663 101 669 106
rect 677 101 693 106
rect 677 88 682 101
rect 668 42 673 48
rect 668 38 682 42
rect 688 41 693 101
rect 709 101 714 115
rect 733 106 736 111
rect 744 106 749 119
rect 773 128 822 131
rect 773 116 778 128
rect 819 125 909 128
rect 796 122 813 125
rect 744 102 756 106
rect 744 101 749 102
rect 709 98 749 101
rect 698 92 701 97
rect 709 88 714 98
rect 721 91 737 95
rect 700 41 705 48
rect 721 41 725 91
rect 744 88 749 98
rect 753 57 756 102
rect 782 70 787 76
rect 796 70 799 122
rect 808 116 813 122
rect 840 116 845 125
rect 872 116 877 125
rect 904 116 909 125
rect 782 67 799 70
rect 807 63 809 68
rect 782 60 803 63
rect 817 60 822 76
rect 849 68 854 76
rect 839 63 841 68
rect 849 63 873 68
rect 881 64 886 76
rect 913 67 918 76
rect 913 64 924 67
rect 849 60 854 63
rect 753 53 774 57
rect 782 50 787 60
rect 800 57 822 60
rect 828 57 854 60
rect 881 59 905 64
rect 735 43 740 48
rect 688 38 725 41
rect 588 34 614 35
rect 460 31 614 34
rect 588 30 614 31
rect 622 32 641 37
rect 309 19 327 23
rect 343 19 359 23
rect 375 19 391 23
rect 460 15 474 18
rect 236 0 241 7
rect 269 3 438 6
rect 236 -4 250 0
rect 159 -24 177 -20
rect 193 -24 209 -20
rect 269 -27 273 3
rect 276 -3 430 0
rect 116 -30 273 -27
rect 282 -9 287 -3
rect 314 -9 319 -3
rect 346 -9 351 -3
rect 378 -9 383 -3
rect 410 -9 415 -3
rect 30 -42 152 -39
rect -155 -54 -143 -49
rect -226 -63 -195 -58
rect -277 -86 -262 -81
rect -214 -82 -209 -63
rect -149 -81 -143 -54
rect -140 -49 -72 -44
rect 36 -48 41 -42
rect 68 -48 73 -42
rect 100 -48 105 -42
rect 132 -48 137 -42
rect 163 -48 166 -43
rect -140 -56 -137 -49
rect -140 -61 -130 -56
rect -86 -57 -81 -54
rect -140 -77 -137 -61
rect -23 -61 -12 -56
rect -90 -70 -63 -65
rect -140 -81 -83 -77
rect -155 -86 -143 -81
rect -222 -95 -195 -90
rect -214 -117 -209 -95
rect -149 -101 -143 -86
rect -135 -96 -130 -91
rect -87 -93 -83 -81
rect -80 -100 -77 -70
rect 434 -26 438 3
rect 433 -29 439 -26
rect 162 -58 252 -52
rect -72 -92 -67 -89
rect -19 -96 -8 -91
rect -90 -105 -59 -100
rect 30 -102 37 -97
rect -77 -111 -72 -105
rect 45 -106 50 -88
rect 66 -102 69 -97
rect 77 -106 82 -88
rect 98 -102 101 -97
rect 109 -106 114 -88
rect 141 -102 146 -88
rect 168 -64 173 -58
rect 200 -64 205 -58
rect 232 -64 237 -58
rect 279 -63 283 -58
rect 126 -106 133 -104
rect 45 -109 133 -106
rect 141 -107 158 -102
rect 291 -66 296 -49
rect 312 -63 315 -58
rect 323 -66 328 -49
rect 344 -63 347 -58
rect 355 -66 360 -49
rect 376 -63 379 -58
rect 387 -65 392 -49
rect 419 -63 424 -49
rect 387 -66 411 -65
rect 291 -69 411 -66
rect 387 -70 411 -69
rect 419 -68 430 -63
rect 291 -79 305 -76
rect 45 -116 59 -112
rect -429 -141 -412 -138
rect -473 -144 -454 -141
rect -537 -148 -532 -145
rect -619 -155 -612 -151
rect -604 -158 -599 -148
rect -586 -151 -564 -148
rect -558 -151 -532 -148
rect -505 -149 -481 -144
rect -594 -154 -589 -152
rect -571 -154 -566 -151
rect -586 -161 -575 -158
rect -558 -156 -554 -151
rect -563 -159 -554 -156
rect -541 -154 -536 -151
rect -518 -154 -513 -152
rect -586 -162 -581 -161
rect -613 -192 -608 -188
rect -578 -192 -575 -161
rect -563 -162 -558 -159
rect -533 -161 -522 -158
rect -505 -156 -500 -149
rect -473 -152 -468 -144
rect -404 -145 -402 -140
rect -429 -148 -408 -145
rect -394 -148 -389 -132
rect -362 -140 -357 -132
rect -372 -145 -370 -140
rect -362 -145 -338 -140
rect -330 -144 -325 -132
rect -298 -141 -293 -132
rect -362 -148 -357 -145
rect -510 -159 -500 -156
rect -533 -162 -528 -161
rect -525 -192 -522 -161
rect -510 -162 -505 -159
rect -443 -155 -437 -151
rect -429 -158 -424 -148
rect -411 -151 -389 -148
rect -383 -151 -357 -148
rect -330 -149 -306 -144
rect -298 -146 -287 -141
rect -613 -195 -590 -192
rect -578 -195 -567 -192
rect -594 -198 -590 -195
rect -542 -198 -537 -192
rect -525 -195 -514 -192
rect -482 -198 -477 -182
rect -419 -154 -414 -152
rect -396 -154 -391 -151
rect -411 -161 -400 -158
rect -383 -156 -379 -151
rect -388 -159 -379 -156
rect -366 -154 -361 -151
rect -343 -154 -338 -152
rect -411 -162 -406 -161
rect -438 -192 -433 -188
rect -403 -192 -400 -161
rect -388 -162 -383 -159
rect -358 -161 -347 -158
rect -330 -156 -325 -149
rect -298 -152 -293 -146
rect -335 -159 -325 -156
rect -358 -162 -353 -161
rect -350 -192 -347 -161
rect -335 -162 -330 -159
rect -277 -150 -263 -145
rect -209 -146 -204 -140
rect -149 -145 -143 -139
rect -438 -195 -415 -192
rect -403 -195 -392 -192
rect -594 -201 -477 -198
rect -419 -198 -415 -195
rect -367 -198 -362 -192
rect -350 -195 -339 -192
rect -307 -198 -302 -182
rect -419 -201 -302 -198
rect -277 -209 -273 -150
rect -155 -150 -143 -145
rect -223 -162 -219 -154
rect -270 -166 -219 -162
rect -209 -159 -195 -154
rect -209 -165 -204 -159
rect -270 -182 -266 -166
rect -215 -170 -204 -165
rect -223 -178 -218 -175
rect -215 -186 -212 -170
rect -209 -178 -204 -175
rect -149 -177 -143 -150
rect -140 -157 -130 -152
rect -77 -153 -72 -147
rect -17 -152 -11 -146
rect -140 -166 -136 -157
rect -23 -157 -11 -152
rect -90 -166 -63 -161
rect -77 -172 -72 -166
rect -17 -172 -11 -157
rect -155 -182 -143 -177
rect -226 -191 -195 -186
rect -277 -214 -262 -209
rect -214 -210 -209 -191
rect -149 -209 -143 -182
rect -140 -177 -72 -172
rect -140 -184 -137 -177
rect 36 -180 41 -176
rect -140 -189 -130 -184
rect -86 -185 -81 -182
rect -140 -205 -137 -189
rect -23 -189 -12 -184
rect 36 -186 50 -180
rect 55 -182 59 -116
rect 66 -119 69 -114
rect 77 -122 93 -118
rect 98 -119 101 -114
rect 109 -122 114 -109
rect 141 -115 146 -107
rect 89 -182 93 -122
rect 132 -162 137 -155
rect 132 -166 146 -162
rect 55 -186 73 -182
rect 89 -186 105 -182
rect -90 -198 -63 -193
rect 30 -195 120 -189
rect 155 -191 158 -107
rect 177 -113 182 -104
rect 166 -118 169 -113
rect 177 -118 193 -113
rect 198 -118 201 -113
rect 209 -118 214 -104
rect 241 -118 246 -104
rect 188 -121 193 -118
rect 209 -121 233 -118
rect 188 -123 233 -121
rect 241 -123 252 -118
rect 188 -124 214 -123
rect 177 -132 189 -128
rect 198 -132 201 -127
rect 168 -182 173 -172
rect 185 -175 189 -132
rect 209 -135 214 -124
rect 241 -131 246 -123
rect 185 -179 205 -175
rect 232 -182 237 -171
rect 168 -186 237 -182
rect 155 -194 234 -191
rect -140 -209 -83 -205
rect -155 -214 -143 -209
rect -222 -223 -195 -218
rect -214 -245 -209 -223
rect -149 -229 -143 -214
rect -135 -224 -130 -219
rect -87 -221 -83 -209
rect -80 -228 -77 -198
rect 36 -201 41 -195
rect 68 -201 73 -195
rect 100 -201 105 -195
rect 149 -200 198 -197
rect -72 -220 -67 -217
rect -19 -224 -8 -219
rect -90 -233 -59 -228
rect -77 -239 -72 -233
rect 149 -203 152 -200
rect 195 -203 198 -200
rect 126 -206 152 -203
rect 155 -206 189 -203
rect 195 -206 221 -203
rect 228 -204 234 -194
rect 45 -250 50 -241
rect 30 -255 37 -250
rect 45 -255 61 -250
rect 66 -255 69 -250
rect 77 -255 82 -241
rect 56 -258 61 -255
rect 77 -258 101 -255
rect 56 -260 101 -258
rect 56 -261 82 -260
rect -177 -264 -128 -261
rect -177 -276 -172 -264
rect -131 -267 -41 -264
rect -154 -270 -137 -267
rect -168 -322 -163 -316
rect -154 -322 -151 -270
rect -142 -276 -137 -270
rect -110 -276 -105 -267
rect -78 -276 -73 -267
rect -46 -276 -41 -267
rect 45 -269 57 -265
rect 66 -269 69 -264
rect -168 -325 -151 -322
rect -143 -329 -141 -324
rect -168 -332 -147 -329
rect -133 -332 -128 -316
rect -101 -324 -96 -316
rect -111 -329 -109 -324
rect -101 -329 -77 -324
rect -69 -328 -64 -316
rect -37 -325 -32 -316
rect 36 -319 41 -309
rect 53 -312 57 -269
rect 77 -272 82 -261
rect 109 -261 114 -241
rect 132 -212 137 -206
rect 141 -261 146 -252
rect 155 -261 160 -206
rect 169 -212 174 -206
rect 201 -212 206 -206
rect 178 -260 183 -252
rect 109 -266 133 -261
rect 141 -266 160 -261
rect 163 -266 170 -261
rect 178 -264 192 -260
rect 188 -266 192 -264
rect 210 -266 215 -252
rect 249 -255 252 -123
rect 282 -163 287 -159
rect 282 -169 296 -163
rect 301 -165 305 -79
rect 312 -82 315 -77
rect 323 -85 339 -81
rect 344 -82 347 -77
rect 355 -85 371 -81
rect 376 -82 379 -77
rect 387 -85 392 -70
rect 419 -78 424 -68
rect 335 -165 339 -85
rect 367 -165 371 -85
rect 410 -122 415 -118
rect 410 -125 424 -122
rect 427 -128 430 -68
rect 451 -89 456 -85
rect 451 -95 465 -89
rect 470 -91 474 15
rect 481 12 484 17
rect 492 9 508 13
rect 513 12 516 17
rect 524 9 540 13
rect 545 12 548 17
rect 556 9 572 13
rect 577 12 580 17
rect 588 9 593 30
rect 622 16 627 32
rect 662 16 688 22
rect 504 -91 508 9
rect 536 -91 540 9
rect 470 -95 488 -91
rect 504 -95 520 -91
rect 536 -95 552 -91
rect 568 -92 572 9
rect 668 10 673 16
rect 700 10 705 21
rect 735 14 740 25
rect 792 54 797 56
rect 815 54 820 57
rect 800 47 811 50
rect 828 52 832 57
rect 823 49 832 52
rect 845 54 850 57
rect 868 54 873 56
rect 800 46 805 47
rect 773 16 778 20
rect 808 16 811 47
rect 823 46 828 49
rect 853 47 864 50
rect 881 52 886 59
rect 913 56 918 64
rect 876 49 886 52
rect 853 46 858 47
rect 861 16 864 47
rect 876 46 881 49
rect 613 -30 618 -24
rect 773 13 796 16
rect 808 13 819 16
rect 792 10 796 13
rect 844 10 849 16
rect 861 13 872 16
rect 904 10 909 26
rect 792 7 909 10
rect 599 -35 618 -30
rect 579 -92 584 -91
rect 568 -95 584 -92
rect 461 -98 465 -95
rect 599 -98 602 -35
rect 677 -39 682 -30
rect 663 -44 669 -39
rect 677 -44 693 -39
rect 677 -57 682 -44
rect 461 -101 602 -98
rect 668 -103 673 -97
rect 668 -107 682 -103
rect 688 -104 693 -44
rect 709 -44 714 -30
rect 733 -39 736 -34
rect 744 -39 749 -26
rect 773 -3 822 0
rect 773 -15 778 -3
rect 819 -6 909 -3
rect 796 -9 813 -6
rect 744 -42 756 -39
rect 744 -44 749 -42
rect 709 -47 749 -44
rect 698 -53 701 -48
rect 709 -57 714 -47
rect 721 -54 737 -50
rect 700 -104 705 -97
rect 721 -104 725 -54
rect 744 -57 749 -47
rect 753 -74 756 -42
rect 782 -61 787 -55
rect 796 -61 799 -9
rect 808 -15 813 -9
rect 840 -15 845 -6
rect 872 -15 877 -6
rect 904 -15 909 -6
rect 782 -64 799 -61
rect 807 -68 809 -63
rect 782 -71 803 -68
rect 817 -71 822 -55
rect 849 -63 854 -55
rect 839 -68 841 -63
rect 849 -68 873 -63
rect 881 -67 886 -55
rect 913 -64 918 -55
rect 913 -67 924 -64
rect 849 -71 854 -68
rect 753 -78 774 -74
rect 782 -81 787 -71
rect 800 -74 822 -71
rect 828 -74 854 -71
rect 881 -72 905 -67
rect 735 -102 740 -97
rect 688 -107 725 -104
rect 792 -77 797 -75
rect 815 -77 820 -74
rect 800 -84 811 -81
rect 828 -79 832 -74
rect 823 -82 832 -79
rect 845 -77 850 -74
rect 868 -77 873 -75
rect 800 -85 805 -84
rect 773 -115 778 -111
rect 808 -115 811 -84
rect 823 -85 828 -82
rect 853 -84 864 -81
rect 881 -79 886 -72
rect 913 -75 918 -67
rect 876 -82 886 -79
rect 853 -85 858 -84
rect 861 -115 864 -84
rect 876 -85 881 -82
rect 773 -118 796 -115
rect 808 -118 819 -115
rect 792 -121 796 -118
rect 844 -121 849 -115
rect 861 -118 872 -115
rect 904 -121 909 -105
rect 403 -131 430 -128
rect 639 -131 665 -125
rect 301 -169 319 -165
rect 335 -169 351 -165
rect 367 -169 383 -165
rect 265 -177 291 -174
rect 294 -177 326 -174
rect 329 -177 361 -174
rect 271 -183 276 -177
rect 280 -253 285 -243
rect 294 -253 297 -177
rect 306 -183 311 -177
rect 249 -260 272 -255
rect 280 -256 297 -253
rect 304 -257 307 -252
rect 315 -253 320 -243
rect 329 -253 332 -177
rect 341 -183 346 -177
rect 367 -204 393 -201
rect 315 -256 332 -253
rect 339 -257 342 -252
rect 350 -262 355 -243
rect 373 -210 378 -204
rect 280 -265 355 -262
rect 109 -268 114 -266
rect 188 -271 202 -266
rect 210 -271 221 -266
rect 188 -274 192 -271
rect 141 -279 154 -276
rect 178 -278 192 -274
rect 141 -280 157 -279
rect 178 -280 183 -278
rect 210 -279 215 -271
rect 280 -276 285 -265
rect 304 -274 307 -269
rect 53 -316 73 -312
rect 100 -319 105 -308
rect 36 -323 105 -319
rect 149 -284 157 -280
rect 315 -277 320 -265
rect 350 -266 355 -265
rect 382 -264 387 -250
rect 403 -260 406 -131
rect 645 -137 650 -131
rect 677 -137 682 -126
rect 712 -133 717 -122
rect 792 -124 909 -121
rect 427 -143 453 -140
rect 456 -143 488 -140
rect 491 -143 523 -140
rect 526 -143 558 -140
rect 433 -149 438 -143
rect 442 -239 447 -229
rect 456 -239 459 -143
rect 468 -149 473 -143
rect 416 -246 434 -241
rect 442 -242 459 -239
rect 466 -243 469 -238
rect 477 -239 482 -229
rect 491 -239 494 -143
rect 503 -149 508 -143
rect 477 -242 494 -239
rect 501 -243 504 -238
rect 512 -239 517 -229
rect 526 -239 529 -143
rect 538 -149 543 -143
rect 654 -186 659 -177
rect 564 -190 590 -187
rect 512 -242 529 -239
rect 533 -243 539 -238
rect 547 -247 552 -229
rect 570 -196 575 -190
rect 640 -191 646 -186
rect 654 -191 670 -186
rect 654 -204 659 -191
rect 547 -248 571 -247
rect 442 -251 571 -248
rect 339 -274 342 -269
rect 350 -271 374 -266
rect 382 -269 390 -264
rect 442 -266 447 -251
rect 466 -264 469 -259
rect 350 -277 355 -271
rect 382 -277 387 -269
rect -37 -328 -18 -325
rect -101 -332 -96 -329
rect -183 -339 -176 -335
rect -168 -342 -163 -332
rect -150 -335 -128 -332
rect -122 -335 -96 -332
rect -69 -333 -45 -328
rect -158 -338 -153 -336
rect -135 -338 -130 -335
rect -150 -345 -139 -342
rect -122 -340 -118 -335
rect -127 -343 -118 -340
rect -105 -338 -100 -335
rect -82 -338 -77 -336
rect -150 -346 -145 -345
rect -177 -376 -172 -372
rect -142 -376 -139 -345
rect -127 -346 -122 -343
rect -97 -345 -86 -342
rect -69 -340 -64 -333
rect -37 -336 -32 -328
rect -24 -333 -18 -328
rect 132 -326 137 -320
rect 169 -326 174 -320
rect 201 -326 206 -319
rect 271 -321 276 -316
rect 477 -267 482 -251
rect 501 -264 504 -259
rect 512 -267 517 -251
rect 547 -252 571 -251
rect 579 -250 584 -236
rect 645 -250 650 -244
rect 533 -264 539 -259
rect 547 -267 552 -252
rect 579 -255 590 -250
rect 645 -254 659 -250
rect 665 -251 670 -191
rect 686 -191 691 -177
rect 710 -186 713 -181
rect 721 -186 726 -173
rect 773 -135 822 -132
rect 773 -147 778 -135
rect 819 -138 909 -135
rect 796 -141 813 -138
rect 721 -191 738 -186
rect 686 -194 726 -191
rect 675 -200 678 -195
rect 686 -204 691 -194
rect 698 -201 714 -197
rect 677 -251 682 -244
rect 698 -251 702 -201
rect 721 -204 726 -194
rect 732 -206 738 -191
rect 782 -193 787 -187
rect 796 -193 799 -141
rect 808 -147 813 -141
rect 840 -147 845 -138
rect 872 -147 877 -138
rect 904 -147 909 -138
rect 782 -196 799 -193
rect 807 -200 809 -195
rect 782 -203 803 -200
rect 817 -203 822 -187
rect 849 -195 854 -187
rect 839 -200 841 -195
rect 849 -200 873 -195
rect 881 -199 886 -187
rect 913 -196 918 -187
rect 913 -199 924 -196
rect 849 -203 854 -200
rect 732 -210 774 -206
rect 782 -213 787 -203
rect 800 -206 822 -203
rect 828 -206 854 -203
rect 881 -204 905 -199
rect 792 -209 797 -207
rect 815 -209 820 -206
rect 800 -216 811 -213
rect 828 -211 832 -206
rect 823 -214 832 -211
rect 845 -209 850 -206
rect 868 -209 873 -207
rect 800 -217 805 -216
rect 712 -249 717 -244
rect 773 -247 778 -243
rect 808 -247 811 -216
rect 823 -217 828 -214
rect 853 -216 864 -213
rect 881 -211 886 -204
rect 913 -207 918 -199
rect 876 -214 886 -211
rect 853 -217 858 -216
rect 861 -247 864 -216
rect 876 -217 881 -214
rect 773 -250 796 -247
rect 808 -250 819 -247
rect 665 -254 702 -251
rect 792 -253 796 -250
rect 844 -253 849 -247
rect 861 -250 872 -247
rect 904 -253 909 -237
rect 579 -267 584 -255
rect 792 -256 909 -253
rect 773 -266 822 -263
rect 433 -311 438 -306
rect 639 -276 665 -270
rect 645 -282 650 -276
rect 677 -282 682 -271
rect 712 -278 717 -267
rect 773 -278 778 -266
rect 819 -269 909 -266
rect 796 -272 813 -269
rect 468 -311 473 -307
rect 503 -311 508 -307
rect 538 -311 543 -307
rect 570 -311 575 -307
rect 433 -314 575 -311
rect 306 -321 311 -317
rect 341 -321 346 -317
rect 373 -321 378 -317
rect 271 -324 378 -321
rect 132 -329 206 -326
rect 654 -331 659 -322
rect 640 -336 646 -331
rect 654 -336 670 -331
rect -74 -343 -64 -340
rect -97 -346 -92 -345
rect -89 -376 -86 -345
rect -74 -346 -69 -343
rect 654 -349 659 -336
rect -177 -379 -154 -376
rect -142 -379 -131 -376
rect -158 -382 -154 -379
rect -106 -382 -101 -376
rect -89 -379 -78 -376
rect -46 -382 -41 -366
rect -158 -385 -41 -382
rect 645 -395 650 -389
rect 645 -399 659 -395
rect 665 -396 670 -336
rect 686 -336 691 -322
rect 710 -331 713 -326
rect 721 -331 726 -318
rect 782 -324 787 -318
rect 796 -324 799 -272
rect 808 -278 813 -272
rect 840 -278 845 -269
rect 872 -278 877 -269
rect 904 -278 909 -269
rect 782 -327 799 -324
rect 807 -331 809 -326
rect 721 -336 738 -331
rect 686 -339 726 -336
rect 675 -345 678 -340
rect 686 -349 691 -339
rect 698 -346 714 -342
rect 677 -396 682 -389
rect 698 -396 702 -346
rect 721 -349 726 -339
rect 732 -337 738 -336
rect 782 -334 803 -331
rect 817 -334 822 -318
rect 849 -326 854 -318
rect 839 -331 841 -326
rect 849 -331 873 -326
rect 881 -330 886 -318
rect 913 -327 918 -318
rect 913 -330 924 -327
rect 849 -334 854 -331
rect 732 -341 774 -337
rect 782 -344 787 -334
rect 800 -337 822 -334
rect 828 -337 854 -334
rect 881 -335 905 -330
rect 792 -340 797 -338
rect 815 -340 820 -337
rect 800 -347 811 -344
rect 828 -342 832 -337
rect 823 -345 832 -342
rect 845 -340 850 -337
rect 868 -340 873 -338
rect 800 -348 805 -347
rect 773 -378 778 -374
rect 808 -378 811 -347
rect 823 -348 828 -345
rect 853 -347 864 -344
rect 881 -342 886 -335
rect 913 -338 918 -330
rect 876 -345 886 -342
rect 853 -348 858 -347
rect 861 -378 864 -347
rect 876 -348 881 -345
rect 773 -381 796 -378
rect 808 -381 819 -378
rect 792 -384 796 -381
rect 844 -384 849 -378
rect 861 -381 872 -378
rect 904 -384 909 -368
rect 792 -387 909 -384
rect 712 -394 717 -389
rect 665 -399 702 -396
<< metal2 >>
rect -459 257 -274 260
rect -459 253 -454 257
rect -277 253 -274 257
rect -277 250 -72 253
rect -209 241 -204 250
rect -77 245 -72 250
rect -77 241 -5 245
rect -77 234 -72 241
rect -9 200 -5 241
rect 196 212 199 222
rect 127 209 199 212
rect 196 200 199 209
rect 421 202 427 205
rect 421 200 451 202
rect -12 195 -5 200
rect 424 199 451 200
rect -9 179 -5 195
rect -72 176 -5 179
rect 448 176 451 199
rect 529 176 532 189
rect -72 167 -67 176
rect 448 173 532 176
rect 529 159 532 173
rect 656 169 724 173
rect -459 127 -274 130
rect -459 122 -454 127
rect -277 125 -274 127
rect 346 125 352 130
rect -277 122 -72 125
rect -209 113 -204 122
rect -77 117 -72 122
rect 346 120 349 125
rect 269 117 349 120
rect -77 113 -5 117
rect -77 106 -72 113
rect -9 72 -5 113
rect -12 67 -5 72
rect -9 51 -5 67
rect 199 55 202 65
rect 120 52 202 55
rect -72 48 -5 51
rect -72 39 -67 48
rect 199 43 202 52
rect 269 5 274 117
rect 346 111 349 117
rect 656 114 659 169
rect 700 166 705 169
rect 346 106 352 111
rect 651 109 659 114
rect 656 106 659 109
rect 721 111 724 169
rect 721 106 733 111
rect 656 101 666 106
rect 507 37 513 42
rect 507 32 510 37
rect 406 29 510 32
rect 406 5 409 29
rect 507 17 510 29
rect 656 24 724 28
rect 531 18 563 21
rect 507 12 513 17
rect 531 16 534 18
rect 560 16 563 18
rect 269 1 409 5
rect -459 -6 -72 -3
rect -459 -10 -454 -6
rect -209 -15 -204 -6
rect -77 -11 -72 -6
rect -77 -15 -5 -11
rect -77 -22 -72 -15
rect -9 -56 -5 -15
rect -12 -61 -5 -56
rect -9 -77 -5 -61
rect 269 -68 274 1
rect 433 -32 439 -29
rect 656 -31 659 24
rect 700 21 705 24
rect 338 -63 344 -58
rect 338 -68 341 -63
rect 269 -71 341 -68
rect 269 -76 274 -71
rect -72 -80 -5 -77
rect 266 -79 274 -76
rect -72 -89 -67 -80
rect 95 -107 98 -97
rect 30 -110 98 -107
rect 30 -112 35 -110
rect 95 -119 98 -110
rect -459 -134 -72 -131
rect -459 -141 -454 -134
rect -209 -143 -204 -134
rect -77 -139 -72 -134
rect -77 -143 -5 -139
rect -77 -150 -72 -143
rect -9 -184 -5 -143
rect 269 -165 274 -79
rect 338 -77 341 -71
rect 338 -82 344 -77
rect 434 -130 438 -32
rect 651 -36 659 -31
rect 656 -39 659 -36
rect 721 -34 724 24
rect 721 -39 733 -34
rect 656 -44 666 -39
rect 407 -133 438 -130
rect 633 -123 701 -119
rect -12 -189 -5 -184
rect -9 -205 -5 -189
rect -72 -208 -5 -205
rect -72 -217 -67 -208
rect 180 -268 188 -266
rect 163 -271 188 -268
rect 228 -270 234 -204
rect 407 -251 410 -133
rect 633 -178 636 -123
rect 677 -126 682 -123
rect 629 -183 636 -178
rect 633 -186 636 -183
rect 698 -181 701 -123
rect 698 -186 710 -181
rect 633 -191 643 -186
rect 498 -251 501 -238
rect 336 -265 339 -252
rect 407 -254 501 -251
rect 498 -264 501 -254
rect 265 -268 339 -265
rect 265 -270 269 -268
rect 163 -272 184 -271
rect 163 -279 166 -272
rect 228 -276 269 -270
rect 336 -274 339 -268
rect 633 -268 701 -264
rect 157 -284 166 -279
rect 633 -323 636 -268
rect 677 -271 682 -268
rect 619 -328 636 -323
rect 633 -331 636 -328
rect 698 -326 701 -268
rect 698 -331 710 -326
rect 633 -336 643 -331
<< metal3 >>
rect -450 318 762 324
rect -585 252 -579 254
rect -623 249 -579 252
rect -553 249 -547 254
rect -450 252 -447 318
rect 6 285 261 288
rect -410 252 -404 254
rect -450 249 -404 252
rect -378 249 -372 254
rect -287 249 -284 251
rect -623 121 -620 249
rect -594 242 -589 249
rect -585 245 -582 249
rect -553 245 -550 249
rect -585 242 -513 245
rect -585 121 -579 123
rect -623 118 -579 121
rect -553 118 -547 123
rect -450 121 -447 249
rect -419 242 -414 249
rect -410 245 -407 249
rect -378 245 -375 249
rect -287 246 -81 249
rect -410 242 -338 245
rect -217 212 -212 246
rect -223 209 -204 212
rect -86 211 -81 246
rect -86 207 0 211
rect -86 202 -81 207
rect -3 175 0 207
rect -83 172 0 175
rect -142 169 -80 172
rect -142 165 -138 169
rect -3 165 0 172
rect -142 160 -135 165
rect -8 160 0 165
rect -410 121 -404 123
rect -450 118 -404 121
rect -378 118 -372 123
rect -287 121 -284 122
rect -287 118 -81 121
rect -623 -11 -620 118
rect -594 111 -589 118
rect -585 114 -582 118
rect -553 114 -550 118
rect -585 111 -513 114
rect -585 -11 -579 -9
rect -623 -14 -579 -11
rect -553 -14 -547 -9
rect -450 -11 -447 118
rect -419 111 -414 118
rect -410 114 -407 118
rect -378 114 -375 118
rect -287 117 -284 118
rect -410 111 -338 114
rect -217 84 -212 118
rect -223 81 -204 84
rect -86 83 -81 118
rect -86 79 0 83
rect -86 74 -81 79
rect -3 47 0 79
rect -83 44 0 47
rect -142 41 -80 44
rect -142 37 -138 41
rect -3 37 0 44
rect -142 32 -135 37
rect -8 32 0 37
rect -410 -11 -404 -9
rect -450 -14 -404 -11
rect -378 -14 -372 -9
rect -278 -10 -81 -7
rect -623 -142 -620 -14
rect -594 -21 -589 -14
rect -585 -18 -582 -14
rect -553 -18 -550 -14
rect -585 -21 -513 -18
rect -585 -142 -579 -140
rect -623 -145 -579 -142
rect -553 -145 -547 -140
rect -450 -142 -447 -14
rect -419 -21 -414 -14
rect -410 -18 -407 -14
rect -378 -18 -375 -14
rect -287 -15 -275 -10
rect -410 -21 -338 -18
rect -217 -44 -212 -10
rect -223 -47 -204 -44
rect -86 -45 -81 -10
rect -86 -49 0 -45
rect -86 -54 -81 -49
rect -3 -81 0 -49
rect -83 -84 0 -81
rect -142 -87 -80 -84
rect -142 -91 -138 -87
rect -3 -91 0 -84
rect -142 -96 -135 -91
rect -8 -96 0 -91
rect 6 -64 12 285
rect 164 216 167 222
rect 123 213 167 216
rect 53 189 56 197
rect 17 184 56 189
rect 17 178 22 184
rect 53 178 56 184
rect 123 136 126 213
rect 164 200 167 213
rect 258 196 261 285
rect 294 240 378 318
rect 756 198 762 318
rect 801 198 807 200
rect 258 193 445 196
rect 442 142 445 193
rect 756 195 807 198
rect 833 195 839 200
rect 756 192 766 195
rect 494 180 497 189
rect 454 177 497 180
rect 454 145 457 177
rect 494 159 497 177
rect 689 175 740 178
rect 110 133 126 136
rect 439 138 445 142
rect 451 142 457 145
rect 110 123 113 133
rect 314 125 320 130
rect 314 124 317 125
rect 21 120 113 123
rect 160 121 317 124
rect 21 41 24 120
rect 160 59 163 121
rect 314 111 317 121
rect 314 106 320 111
rect 167 59 170 65
rect 439 62 442 138
rect 451 131 454 142
rect 449 128 454 131
rect 689 97 693 175
rect 725 98 728 175
rect 735 170 740 175
rect 656 92 698 97
rect 725 95 731 98
rect 656 89 661 92
rect 130 56 170 59
rect 61 41 64 49
rect 21 36 64 41
rect 61 30 64 36
rect 130 -32 134 56
rect 167 43 170 56
rect 435 59 442 62
rect 435 36 438 59
rect 475 37 481 42
rect 728 40 731 95
rect 763 66 766 192
rect 792 188 797 195
rect 801 191 804 195
rect 833 191 836 195
rect 801 188 873 191
rect 801 66 807 68
rect 763 63 807 66
rect 833 63 839 68
rect 735 40 740 43
rect 728 37 740 40
rect 475 36 478 37
rect 435 33 478 36
rect 262 25 267 28
rect 263 10 266 25
rect 475 17 478 33
rect 689 30 740 33
rect 475 12 481 17
rect 263 7 443 10
rect 130 -37 182 -32
rect 179 -43 182 -37
rect 176 -48 182 -43
rect 306 -63 312 -58
rect 306 -64 309 -63
rect 6 -67 309 -64
rect 6 -103 12 -67
rect 306 -77 309 -67
rect 306 -82 312 -77
rect 63 -103 66 -97
rect 6 -106 66 -103
rect -283 -138 -81 -135
rect -410 -142 -404 -140
rect -450 -145 -404 -142
rect -378 -145 -372 -140
rect -283 -141 -280 -138
rect -623 -202 -620 -145
rect -594 -152 -589 -145
rect -585 -149 -582 -145
rect -553 -149 -550 -145
rect -585 -152 -513 -149
rect -450 -202 -447 -145
rect -419 -152 -414 -145
rect -410 -149 -407 -145
rect -378 -149 -375 -145
rect -287 -146 -280 -141
rect -410 -152 -338 -149
rect -217 -172 -212 -138
rect -223 -175 -204 -172
rect -86 -173 -81 -138
rect -86 -177 0 -173
rect -86 -182 -81 -177
rect -623 -204 -447 -202
rect -623 -205 -288 -204
rect -450 -210 -288 -205
rect -3 -209 0 -177
rect -294 -228 -288 -210
rect -83 -212 0 -209
rect -142 -215 -80 -212
rect -142 -219 -138 -215
rect -3 -219 0 -212
rect -142 -224 -135 -219
rect -8 -224 0 -219
rect -294 -234 -222 -228
rect -228 -324 -222 -234
rect 6 -258 12 -106
rect 63 -119 66 -106
rect 195 -123 198 -113
rect 168 -126 198 -123
rect 168 -128 171 -126
rect 195 -132 198 -126
rect 440 -132 443 7
rect 689 -48 693 30
rect 725 -47 728 30
rect 735 25 740 30
rect 661 -53 698 -48
rect 725 -50 731 -47
rect 661 -99 664 -53
rect 411 -135 443 -132
rect 628 -107 664 -99
rect 728 -105 731 -50
rect 763 -65 766 63
rect 792 56 797 63
rect 801 59 804 63
rect 833 59 836 63
rect 801 56 873 59
rect 801 -65 807 -63
rect 763 -68 807 -65
rect 833 -68 839 -63
rect 735 -105 740 -102
rect 411 -247 414 -135
rect 628 -172 632 -107
rect 728 -108 740 -105
rect 615 -176 632 -172
rect 666 -117 717 -114
rect 463 -247 466 -238
rect 411 -250 466 -247
rect 63 -258 66 -250
rect 6 -263 66 -258
rect 301 -261 304 -252
rect -228 -326 -186 -324
rect -149 -326 -143 -324
rect -228 -329 -143 -326
rect -117 -329 -111 -324
rect -228 -330 -186 -329
rect -158 -336 -153 -329
rect -149 -333 -146 -329
rect -117 -333 -114 -329
rect -149 -336 -77 -333
rect -24 -339 -18 -333
rect 6 -339 12 -263
rect 63 -269 66 -263
rect 158 -266 163 -261
rect 261 -264 304 -261
rect 463 -264 466 -250
rect 261 -266 264 -264
rect 158 -268 161 -266
rect 126 -273 161 -268
rect 221 -330 224 -266
rect 301 -274 304 -264
rect 390 -321 393 -264
rect 615 -288 619 -176
rect 666 -195 670 -117
rect 702 -194 705 -117
rect 712 -122 717 -117
rect 595 -294 619 -288
rect 629 -200 675 -195
rect 702 -197 708 -194
rect 595 -321 601 -294
rect 629 -312 632 -200
rect 705 -252 708 -197
rect 763 -197 766 -68
rect 792 -75 797 -68
rect 801 -72 804 -68
rect 833 -72 836 -68
rect 801 -75 873 -72
rect 801 -197 807 -195
rect 763 -200 807 -197
rect 833 -200 839 -195
rect 712 -252 717 -249
rect 705 -255 717 -252
rect 390 -324 601 -321
rect 609 -318 632 -312
rect 666 -262 717 -259
rect 609 -330 615 -318
rect 221 -333 615 -330
rect 666 -339 670 -262
rect 702 -339 705 -262
rect 712 -267 717 -262
rect 763 -328 766 -200
rect 792 -207 797 -200
rect 801 -204 804 -200
rect 833 -204 836 -200
rect 801 -207 873 -204
rect 801 -328 807 -326
rect 763 -331 807 -328
rect 833 -331 839 -326
rect 792 -338 797 -331
rect 801 -335 804 -331
rect 833 -335 836 -331
rect 801 -338 873 -335
rect -24 -344 675 -339
rect 702 -342 708 -339
rect 705 -397 708 -342
rect 712 -397 717 -394
rect 705 -400 717 -397
<< metal4 >>
rect 250 212 269 217
rect 266 202 269 212
rect 415 202 421 205
rect 266 200 421 202
rect 266 199 418 200
rect 564 172 567 189
rect 452 169 567 172
rect 452 166 455 169
rect 449 161 455 166
rect 564 159 567 169
rect 381 116 384 130
rect 260 113 384 116
rect 381 106 384 113
rect 656 86 661 89
rect 542 28 545 42
rect 445 25 545 28
rect 410 18 531 21
rect 410 5 414 18
rect 528 16 531 18
rect 542 12 545 25
rect 574 21 577 42
rect 563 18 577 21
rect 563 16 566 18
rect 574 12 577 18
rect 252 2 414 5
rect 252 -58 255 2
rect 252 -63 279 -58
rect 252 -175 255 -63
rect 373 -72 376 -58
rect 265 -75 376 -72
rect 278 -170 281 -75
rect 373 -82 376 -75
rect 657 -110 660 86
rect 633 -118 660 -110
rect 240 -178 255 -175
rect 240 -278 243 -178
rect 634 -225 637 -118
rect 533 -255 536 -238
rect 634 -250 638 -225
rect 590 -255 638 -250
rect 406 -258 536 -255
rect 406 -260 409 -258
rect 533 -264 536 -258
rect 231 -282 243 -278
rect 231 -324 236 -282
<< metal5 >>
rect 124 281 257 284
rect 124 263 129 281
rect 9 260 129 263
rect 9 197 14 260
rect 124 222 129 260
rect 2 192 23 197
rect -77 142 -72 145
rect 2 142 6 192
rect -77 138 6 142
rect 127 127 132 209
rect 254 192 257 281
rect 272 206 277 215
rect 436 209 439 210
rect 410 206 439 209
rect 272 203 413 206
rect 436 205 439 206
rect 254 189 444 192
rect 254 137 257 189
rect 254 134 283 137
rect 278 130 283 134
rect 120 124 260 127
rect 120 114 124 124
rect 160 123 163 124
rect 13 111 124 114
rect -77 14 -72 17
rect 13 14 17 111
rect 119 110 124 111
rect 257 116 260 124
rect 381 116 384 130
rect 257 113 384 116
rect 119 69 122 110
rect 119 65 124 69
rect -77 10 17 14
rect 120 -35 125 52
rect 257 14 260 113
rect 381 106 384 113
rect 439 103 444 189
rect 599 168 602 189
rect 456 165 602 168
rect 456 115 460 165
rect 599 159 602 165
rect 455 109 461 115
rect 648 103 651 114
rect 439 100 651 103
rect 439 45 444 100
rect 542 28 545 42
rect 402 25 545 28
rect 402 14 405 25
rect 257 10 405 14
rect 542 12 545 25
rect 257 -25 260 10
rect 257 -28 265 -25
rect 24 -38 162 -35
rect 24 -97 27 -38
rect 2 -102 30 -97
rect -77 -114 -72 -111
rect 2 -114 5 -102
rect -77 -118 5 -114
rect -77 -242 -72 -239
rect 25 -242 30 -107
rect 159 -113 162 -38
rect 167 -48 170 -43
rect 262 -72 265 -28
rect 643 -36 651 -31
rect 373 -72 376 -58
rect 262 -75 376 -72
rect 159 -118 166 -113
rect 159 -197 162 -118
rect 269 -169 274 -165
rect 261 -173 274 -169
rect 278 -170 281 -75
rect 373 -82 376 -75
rect 643 -94 648 -36
rect 623 -98 648 -94
rect 623 -167 627 -98
rect 278 -173 399 -170
rect 261 -197 264 -173
rect 159 -200 264 -197
rect -77 -246 30 -242
rect 25 -334 30 -246
rect 231 -334 236 -324
rect 247 -325 253 -200
rect 396 -316 399 -173
rect 611 -171 627 -167
rect 611 -276 615 -171
rect 588 -282 615 -276
rect 620 -183 629 -178
rect 588 -316 594 -282
rect 620 -300 626 -183
rect 396 -320 594 -316
rect 602 -306 626 -300
rect 602 -325 608 -306
rect 247 -329 608 -325
rect 619 -334 625 -328
rect 25 -338 625 -334
<< metal6 >>
rect 0 289 272 294
rect 0 136 5 289
rect 267 223 272 289
rect 267 218 277 223
rect -214 131 5 136
rect 17 120 22 175
rect 114 127 266 132
rect 114 120 119 127
rect 0 115 119 120
rect 0 8 5 115
rect 261 66 266 127
rect 261 61 273 66
rect 268 41 273 61
rect -214 3 5 8
rect 268 36 277 41
rect 28 -29 33 31
rect 272 16 277 36
rect 272 11 449 16
rect 14 -34 261 -29
rect 14 -120 20 -34
rect 152 -43 157 -39
rect 152 -48 173 -43
rect -214 -125 20 -120
rect 152 -123 157 -48
rect 149 -128 165 -123
rect 149 -189 154 -128
rect 121 -194 154 -189
rect -214 -253 18 -248
rect -6 -326 0 -253
rect 121 -268 126 -194
rect 256 -261 261 -34
rect 444 -133 449 11
rect 416 -138 449 -133
rect 416 -246 421 -138
rect 121 -326 126 -273
rect -6 -331 126 -326
<< pad >>
rect -582 249 -577 254
rect -550 249 -545 254
rect -459 250 -454 255
rect -407 249 -402 254
rect -375 249 -370 254
rect -289 246 -284 251
rect -594 240 -589 245
rect -518 240 -513 245
rect -419 240 -414 245
rect -343 240 -338 245
rect -209 238 -204 244
rect -77 231 -72 237
rect -223 206 -218 212
rect -209 206 -204 212
rect -86 199 -81 204
rect -15 195 -9 200
rect -138 160 -132 165
rect -72 164 -67 170
rect -11 160 -5 165
rect -77 142 -72 148
rect -214 136 -209 142
rect 124 217 129 226
rect 164 217 170 222
rect 196 217 202 222
rect 247 212 253 217
rect 127 206 132 212
rect 272 211 277 218
rect 436 205 442 210
rect 164 200 170 205
rect 196 200 202 205
rect 418 200 424 205
rect 20 192 26 197
rect 53 192 59 197
rect 804 195 809 200
rect 836 195 841 200
rect 494 184 500 189
rect 529 184 535 189
rect 564 184 570 189
rect 599 184 605 189
rect 792 186 797 191
rect 868 186 873 191
rect 17 175 22 181
rect 53 178 59 183
rect -582 118 -577 123
rect -550 118 -545 123
rect -459 119 -454 124
rect -407 118 -402 123
rect -375 118 -370 123
rect -289 117 -284 122
rect 446 161 452 166
rect 494 159 500 164
rect 529 159 535 164
rect 564 159 570 164
rect 599 159 605 164
rect 700 163 705 169
rect 735 167 740 173
rect 278 128 283 133
rect -594 109 -589 114
rect -518 109 -513 114
rect -419 109 -414 114
rect -343 109 -338 114
rect -209 110 -204 116
rect -77 103 -72 109
rect -223 78 -218 84
rect -209 78 -204 84
rect -86 71 -81 76
rect -15 67 -9 72
rect -138 32 -132 37
rect -72 36 -67 42
rect -11 32 -5 37
rect -77 14 -72 20
rect -214 8 -209 14
rect 119 62 124 67
rect 317 125 323 130
rect 349 125 355 130
rect 381 125 387 130
rect 449 125 454 131
rect 317 106 323 111
rect 349 106 355 111
rect 381 106 387 111
rect 455 106 461 112
rect 648 109 654 114
rect 730 106 736 111
rect 663 101 669 106
rect 696 92 701 97
rect 656 86 661 92
rect 167 60 173 65
rect 199 60 205 65
rect 804 63 809 68
rect 836 63 841 68
rect 120 49 125 55
rect 14 44 20 49
rect 61 44 67 49
rect 167 43 173 48
rect 199 43 205 48
rect 792 54 797 59
rect 868 54 873 59
rect 439 42 444 48
rect 28 31 33 41
rect 478 37 484 42
rect 510 37 516 42
rect 542 37 548 42
rect 574 37 580 42
rect 735 40 740 46
rect -582 -14 -577 -9
rect -550 -14 -545 -9
rect -459 -13 -454 -8
rect -407 -14 -402 -9
rect -375 -14 -370 -9
rect -290 -15 -284 -10
rect -209 -18 -204 -12
rect -594 -23 -589 -18
rect -518 -23 -513 -18
rect -419 -23 -414 -18
rect -343 -23 -338 -18
rect -77 -25 -72 -19
rect 61 30 67 35
rect 262 25 267 31
rect 478 12 484 17
rect 510 12 516 17
rect 528 16 534 21
rect 542 12 548 17
rect 560 16 566 21
rect 700 18 705 24
rect 735 22 740 28
rect 574 12 580 17
rect 433 -32 439 -26
rect -223 -50 -218 -44
rect -209 -50 -204 -44
rect -86 -57 -81 -52
rect -15 -61 -9 -56
rect -138 -96 -132 -91
rect -72 -92 -67 -86
rect -11 -96 -5 -91
rect -77 -114 -72 -108
rect -214 -120 -209 -114
rect 173 -48 179 -43
rect 27 -102 33 -97
rect 63 -102 69 -97
rect 95 -102 101 -97
rect 25 -112 35 -107
rect 63 -119 69 -114
rect 95 -119 101 -114
rect 163 -118 169 -113
rect 195 -118 201 -113
rect 165 -128 171 -123
rect -582 -145 -577 -140
rect -550 -145 -545 -140
rect -459 -144 -454 -139
rect -407 -145 -402 -140
rect -375 -145 -370 -140
rect -290 -146 -284 -141
rect -209 -146 -204 -140
rect -594 -154 -589 -149
rect -518 -154 -513 -149
rect -419 -154 -414 -149
rect -343 -154 -338 -149
rect -77 -153 -72 -147
rect -223 -178 -218 -172
rect -209 -178 -204 -172
rect -86 -185 -81 -180
rect -15 -189 -9 -184
rect 195 -132 201 -127
rect -138 -224 -132 -219
rect -72 -220 -67 -214
rect -11 -224 -5 -219
rect -77 -242 -72 -236
rect -214 -248 -209 -242
rect -146 -329 -141 -324
rect -114 -329 -109 -324
rect 25 -255 35 -250
rect 63 -255 69 -250
rect 63 -269 69 -264
rect 228 -207 234 -201
rect 276 -63 282 -58
rect 309 -63 315 -58
rect 341 -63 347 -58
rect 373 -63 379 -58
rect 309 -82 315 -77
rect 341 -82 347 -77
rect 373 -82 379 -77
rect 648 -36 654 -31
rect 730 -39 736 -34
rect 663 -44 669 -39
rect 696 -53 701 -48
rect 804 -68 809 -63
rect 836 -68 841 -63
rect 792 -77 797 -72
rect 868 -77 873 -72
rect 735 -105 740 -99
rect 677 -129 682 -123
rect 712 -125 717 -119
rect 269 -168 274 -162
rect 626 -183 632 -178
rect 707 -186 713 -181
rect 640 -191 646 -186
rect 673 -200 678 -195
rect 804 -200 809 -195
rect 836 -200 841 -195
rect 792 -209 797 -204
rect 868 -209 873 -204
rect 421 -246 427 -241
rect 463 -243 469 -238
rect 498 -243 504 -238
rect 533 -243 539 -238
rect 301 -257 307 -252
rect 336 -257 342 -252
rect 587 -255 593 -250
rect 712 -252 717 -246
rect 403 -260 409 -255
rect 163 -266 168 -261
rect 256 -266 264 -261
rect 463 -264 469 -259
rect 498 -264 504 -259
rect 533 -264 539 -259
rect 121 -273 132 -268
rect 184 -271 192 -266
rect 218 -271 224 -266
rect 387 -269 393 -264
rect 301 -274 307 -269
rect 336 -274 342 -269
rect 677 -274 682 -268
rect 712 -270 717 -264
rect 154 -284 160 -279
rect -158 -338 -153 -333
rect -82 -338 -77 -333
rect -24 -336 -18 -330
rect 231 -327 236 -321
rect 619 -334 625 -323
rect 707 -331 713 -326
rect 804 -331 809 -326
rect 836 -331 841 -326
rect 640 -336 646 -331
rect 792 -340 797 -335
rect 868 -340 873 -335
rect 673 -345 678 -340
rect 712 -397 717 -391
<< labels >>
rlabel metal1 353 -2 353 -2 1 vdd!
rlabel metal1 289 -166 289 -166 1 gnd!
rlabel metal1 417 -124 417 -124 1 gnd!
rlabel metal5 -19 -116 -19 -116 1 p1
rlabel metal6 -19 5 -19 5 1 g2
rlabel metal1 73 -22 73 -22 1 gnd!
rlabel metal1 73 107 73 107 1 vdd!
rlabel metal1 329 -323 329 -323 1 gnd!
rlabel metal1 -146 -184 -146 -184 1 vdd!
rlabel metal1 -146 -56 -146 -56 1 vdd!
rlabel metal1 -146 72 -146 72 1 vdd!
rlabel metal1 -146 200 -146 200 1 vdd!
rlabel metal1 -14 225 -14 225 1 vdd!
rlabel metal1 -14 97 -14 97 1 vdd!
rlabel metal1 -14 -31 -14 -31 1 vdd!
rlabel metal1 -138 -159 -138 -159 1 gnd!
rlabel metal1 -275 -184 -275 -184 3 gnd!
rlabel metal1 -275 -56 -275 -56 3 gnd!
rlabel metal1 -138 -32 -138 -32 1 gnd!
rlabel metal1 -138 97 -138 97 1 gnd!
rlabel metal1 -275 72 -275 72 3 gnd!
rlabel metal1 -275 200 -275 200 3 gnd!
rlabel metal1 -138 225 -138 225 1 gnd!
rlabel metal5 -19 12 -19 12 1 p2
rlabel metal1 195 121 195 121 1 vdd!
rlabel metal1 147 -20 147 -20 1 gnd!
rlabel metal1 243 -2 243 -2 1 gnd!
rlabel metal1 207 -184 207 -184 1 gnd!
rlabel metal1 -14 -159 -14 -159 1 vdd!
rlabel metal1 171 -327 171 -327 1 gnd!
rlabel metal1 75 -321 75 -321 1 gnd!
rlabel metal1 43 -183 43 -183 1 gnd!
rlabel metal1 75 -192 75 -192 1 vdd!
rlabel metal3 -273 -136 -273 -136 3 b0
rlabel metal3 -273 -8 -273 -8 3 b1
rlabel metal2 -273 -5 -273 -5 3 a1
rlabel metal3 -273 120 -273 120 3 b2
rlabel metal2 -273 123 -273 123 3 a2
rlabel metal3 -273 248 -273 248 4 b3
rlabel metal1 440 -142 440 -142 1 vdd!
rlabel metal1 577 -189 577 -189 1 vdd!
rlabel metal1 510 -313 510 -313 1 gnd!
rlabel metal1 652 -273 652 -273 1 vdd!
rlabel metal1 652 -128 652 -128 1 vdd!
rlabel metal1 652 -252 652 -252 1 gnd!
rlabel metal1 652 -397 652 -397 1 gnd!
rlabel metal1 675 164 675 164 1 vdd!
rlabel metal1 675 -105 675 -105 1 gnd!
rlabel metal1 675 40 675 40 1 gnd!
rlabel metal1 675 19 675 19 1 vdd!
rlabel metal1 361 186 361 186 1 vdd!
rlabel metal1 297 22 297 22 1 gnd!
rlabel metal1 425 60 425 60 1 gnd!
rlabel metal1 144 136 144 136 1 gnd!
rlabel metal1 240 155 240 155 1 gnd!
rlabel metal1 65 126 65 126 1 gnd!
rlabel metal1 65 255 65 255 1 vdd!
rlabel metal1 192 279 192 279 5 vdd!
rlabel metal1 154 -199 154 -199 1 vdd!
rlabel metal3 9 -341 9 -341 1 c0
rlabel metal3 223 -331 223 -331 1 c1
rlabel metal3 392 -322 392 -322 1 c2
rlabel metal4 636 -253 636 -253 1 c3
rlabel metal5 -19 140 -19 140 1 p3
rlabel metal6 -19 -122 -19 -122 1 g1
rlabel metal6 -19 -251 -19 -251 1 g0
rlabel metal5 -19 -244 -19 -244 1 p0
rlabel metal1 454 -92 454 -92 1 gnd!
rlabel metal1 538 98 538 98 1 vdd!
rlabel metal1 278 -176 278 -176 1 vdd!
rlabel metal1 541 111 541 111 1 gnd!
rlabel metal1 643 236 643 236 1 vdd!
rlabel metal1 380 -203 380 -203 1 vdd!
rlabel metal1 91 -41 91 -41 1 vdd!
rlabel metal1 208 -55 208 -55 1 vdd!
rlabel metal1 139 -164 139 -164 1 gnd!
rlabel metal6 -19 133 -19 133 1 g3
rlabel metal1 471 405 471 405 5 vdd!
rlabel metal1 -436 201 -436 201 1 gnd!
rlabel metal1 -436 315 -436 315 5 vdd!
rlabel metal1 -414 282 -414 282 1 x1
rlabel metal1 -436 70 -436 70 1 gnd!
rlabel metal1 -436 184 -436 184 5 vdd!
rlabel metal1 -414 151 -414 151 1 x1
rlabel metal1 -414 -112 -414 -112 1 x1
rlabel metal1 -436 -79 -436 -79 5 vdd!
rlabel metal1 -436 -193 -436 -193 1 gnd!
rlabel metal1 -414 19 -414 19 1 x1
rlabel metal1 -436 52 -436 52 5 vdd!
rlabel metal1 -436 -62 -436 -62 1 gnd!
rlabel metal1 -611 201 -611 201 1 gnd!
rlabel metal1 -611 315 -611 315 5 vdd!
rlabel metal1 -589 282 -589 282 1 x1
rlabel metal1 -611 70 -611 70 1 gnd!
rlabel metal1 -611 184 -611 184 5 vdd!
rlabel metal1 -589 151 -589 151 1 x1
rlabel metal1 -589 -112 -589 -112 1 x1
rlabel metal1 -611 -79 -611 -79 5 vdd!
rlabel metal1 -611 -193 -611 -193 1 gnd!
rlabel metal1 -589 19 -589 19 1 x1
rlabel metal1 -611 52 -611 52 5 vdd!
rlabel metal1 -611 -62 -611 -62 1 gnd!
rlabel metal2 -273 -133 -273 -133 3 a0
rlabel metal2 -273 251 -273 251 4 a3
rlabel metal1 -617 241 -617 241 1 a3_in
rlabel metal1 -618 110 -618 110 3 a2_in
rlabel metal1 -618 -22 -618 -22 3 a1_in
rlabel metal1 -618 -153 -618 -153 3 a0_in
rlabel metal1 -442 241 -442 241 1 b3_in
rlabel metal1 -442 110 -442 110 1 b2_in
rlabel metal1 -442 -22 -442 -22 1 b1_in
rlabel metal1 -442 -153 -442 -153 1 b0_in
rlabel metal1 775 15 775 15 1 gnd!
rlabel metal1 775 129 775 129 5 vdd!
rlabel metal1 797 96 797 96 1 x1
rlabel metal1 775 -116 775 -116 1 gnd!
rlabel metal1 775 -2 775 -2 5 vdd!
rlabel metal1 797 -35 797 -35 1 x1
rlabel metal1 797 -298 797 -298 1 x1
rlabel metal1 775 -265 775 -265 5 vdd!
rlabel metal1 775 -379 775 -379 1 gnd!
rlabel metal1 797 -167 797 -167 1 x1
rlabel metal1 775 -134 775 -134 5 vdd!
rlabel metal1 775 -248 775 -248 1 gnd!
rlabel metal1 775 147 775 147 1 gnd!
rlabel metal1 775 261 775 261 5 vdd!
rlabel metal1 797 228 797 228 1 x1
rlabel metal3 336 282 336 282 1 clk
rlabel metal1 921 -329 921 -329 7 s0
rlabel metal1 922 -198 922 -198 7 s1
rlabel metal1 922 -66 922 -66 7 s2
rlabel metal1 922 65 922 65 7 s3
rlabel metal1 922 197 922 197 7 Cout
rlabel metal1 -153 -296 -153 -296 1 x1
rlabel metal1 -175 -263 -175 -263 5 vdd!
rlabel metal1 -175 -377 -175 -377 1 gnd!
rlabel metal1 -182 -337 -182 -337 1 Cin
<< end >>
