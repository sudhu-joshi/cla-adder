magic
tech scmos
timestamp 1733145755
<< nwell >>
rect 312 -202 338 -150
rect 347 -202 373 -150
rect 379 -202 405 -150
rect 411 -202 437 -150
rect 443 -202 469 -150
<< ntransistor >>
rect 324 -252 326 -222
rect 342 -256 344 -226
rect 365 -256 367 -226
rect 395 -256 397 -226
rect 418 -256 420 -226
rect 455 -246 457 -216
<< ptransistor >>
rect 324 -196 326 -156
rect 359 -196 361 -156
rect 391 -196 393 -156
rect 423 -196 425 -156
rect 455 -196 457 -156
<< ndiffusion >>
rect 323 -252 324 -222
rect 326 -252 327 -222
rect 341 -256 342 -226
rect 344 -256 345 -226
rect 364 -256 365 -226
rect 367 -256 368 -226
rect 394 -256 395 -226
rect 397 -256 398 -226
rect 417 -256 418 -226
rect 420 -256 421 -226
rect 454 -246 455 -216
rect 457 -246 458 -216
<< pdiffusion >>
rect 323 -196 324 -156
rect 326 -196 327 -156
rect 358 -196 359 -156
rect 361 -196 362 -156
rect 390 -196 391 -156
rect 393 -196 394 -156
rect 422 -196 423 -156
rect 425 -196 426 -156
rect 454 -196 455 -156
rect 457 -196 458 -156
<< ndcontact >>
rect 318 -252 323 -222
rect 327 -252 332 -222
rect 336 -256 341 -226
rect 345 -256 350 -226
rect 359 -256 364 -226
rect 368 -256 373 -226
rect 389 -256 394 -226
rect 398 -256 403 -226
rect 412 -256 417 -226
rect 421 -256 426 -226
rect 449 -246 454 -216
rect 458 -246 463 -216
<< pdcontact >>
rect 318 -196 323 -156
rect 327 -196 332 -156
rect 353 -196 358 -156
rect 362 -196 367 -156
rect 385 -196 390 -156
rect 394 -196 399 -156
rect 417 -196 422 -156
rect 426 -196 431 -156
rect 449 -196 454 -156
rect 458 -196 463 -156
<< polysilicon >>
rect 324 -156 326 -152
rect 359 -156 361 -152
rect 391 -156 393 -152
rect 423 -156 425 -152
rect 455 -156 457 -152
rect 324 -222 326 -196
rect 359 -209 361 -196
rect 391 -209 393 -196
rect 423 -209 425 -196
rect 455 -216 457 -196
rect 342 -226 344 -218
rect 365 -226 367 -218
rect 395 -226 397 -218
rect 418 -226 420 -218
rect 324 -255 326 -252
rect 455 -249 457 -246
rect 342 -259 344 -256
rect 365 -259 367 -256
rect 395 -259 397 -256
rect 418 -259 420 -256
<< polycontact >>
rect 319 -219 324 -215
rect 354 -209 359 -204
rect 386 -209 391 -204
rect 418 -209 423 -204
rect 450 -213 455 -208
rect 337 -223 342 -218
rect 360 -223 365 -218
rect 390 -223 395 -218
rect 413 -223 418 -218
<< metal1 >>
rect 318 -144 367 -141
rect 318 -156 323 -144
rect 364 -147 454 -144
rect 341 -150 358 -147
rect 327 -202 332 -196
rect 341 -202 344 -150
rect 353 -156 358 -150
rect 385 -156 390 -147
rect 417 -156 422 -147
rect 449 -156 454 -147
rect 327 -205 344 -202
rect 352 -209 354 -204
rect 327 -212 348 -209
rect 362 -212 367 -196
rect 394 -204 399 -196
rect 384 -209 386 -204
rect 394 -209 418 -204
rect 426 -208 431 -196
rect 458 -205 463 -196
rect 458 -208 469 -205
rect 394 -212 399 -209
rect 312 -219 319 -215
rect 327 -222 332 -212
rect 345 -215 367 -212
rect 373 -215 399 -212
rect 426 -213 450 -208
rect 337 -218 342 -216
rect 360 -218 365 -215
rect 345 -225 356 -222
rect 373 -220 377 -215
rect 368 -223 377 -220
rect 390 -218 395 -215
rect 413 -218 418 -216
rect 345 -226 350 -225
rect 318 -256 323 -252
rect 353 -256 356 -225
rect 368 -226 373 -223
rect 398 -225 409 -222
rect 426 -220 431 -213
rect 458 -216 463 -208
rect 421 -223 431 -220
rect 398 -226 403 -225
rect 406 -256 409 -225
rect 421 -226 426 -223
rect 318 -259 341 -256
rect 353 -259 364 -256
rect 337 -262 341 -259
rect 389 -262 394 -256
rect 406 -259 417 -256
rect 449 -262 454 -246
rect 337 -265 454 -262
<< metal3 >>
rect 346 -206 352 -204
rect 312 -209 352 -206
rect 378 -209 384 -204
rect 337 -216 342 -209
rect 346 -213 349 -209
rect 378 -213 381 -209
rect 346 -216 418 -213
<< pad >>
rect 349 -209 354 -204
rect 381 -209 386 -204
rect 337 -218 342 -213
rect 413 -218 418 -213
<< labels >>
rlabel metal1 342 -176 342 -176 1 x1
rlabel metal1 466 -206 466 -206 1 out
rlabel metal1 365 -206 365 -206 1 y1
rlabel metal3 315 -208 315 -208 3 clk
rlabel metal1 320 -143 320 -143 5 vdd!
rlabel metal1 370 -221 370 -221 1 y2
rlabel metal1 320 -257 320 -257 1 gnd!
rlabel metal1 423 -221 423 -221 1 y3
rlabel metal1 354 -242 354 -242 1 x2
rlabel metal1 407 -242 407 -242 1 x3
rlabel metal1 313 -217 313 -217 3 A
<< end >>
