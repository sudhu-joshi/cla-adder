magic
tech scmos
timestamp 1732037377
<< nwell >>
rect -1 30 25 102
rect 34 30 60 102
rect 69 30 95 102
rect 101 23 127 75
<< ntransistor >>
rect 11 -37 13 3
rect 46 -38 48 2
rect 81 -38 83 2
rect 113 -38 115 2
<< ptransistor >>
rect 11 36 13 96
rect 46 36 48 96
rect 81 36 83 96
rect 113 29 115 69
<< ndiffusion >>
rect 10 -37 11 3
rect 13 -37 14 3
rect 45 -38 46 2
rect 48 -38 49 2
rect 80 -38 81 2
rect 83 -38 84 2
rect 112 -38 113 2
rect 115 -38 116 2
<< pdiffusion >>
rect 10 36 11 96
rect 13 36 14 96
rect 45 36 46 96
rect 48 36 49 96
rect 80 36 81 96
rect 83 36 84 96
rect 112 29 113 69
rect 115 29 116 69
<< ndcontact >>
rect 5 -37 10 3
rect 14 -37 19 3
rect 40 -38 45 2
rect 49 -38 54 2
rect 75 -38 80 2
rect 84 -38 89 2
rect 107 -38 112 2
rect 116 -38 121 2
<< pdcontact >>
rect 5 36 10 96
rect 14 36 19 96
rect 40 36 45 96
rect 49 36 54 96
rect 75 36 80 96
rect 84 36 89 96
rect 107 29 112 69
rect 116 29 121 69
<< polysilicon >>
rect 11 96 13 100
rect 46 96 48 100
rect 81 96 83 100
rect 113 69 115 73
rect 11 3 13 36
rect 46 22 48 36
rect 81 22 83 36
rect 46 2 48 10
rect 81 2 83 10
rect 113 2 115 29
rect 11 -40 13 -37
rect 46 -41 48 -38
rect 81 -41 83 -38
rect 113 -41 115 -38
<< polycontact >>
rect 6 19 11 24
rect 41 22 46 27
rect 76 22 81 27
rect 41 5 46 10
rect 76 5 81 10
rect 108 8 113 13
<< metal1 >>
rect -1 102 25 105
rect 28 102 60 105
rect 63 102 95 105
rect 5 96 10 102
rect 14 26 19 36
rect 28 26 31 102
rect 40 96 45 102
rect -1 19 6 24
rect 14 23 31 26
rect 38 22 41 27
rect 49 26 54 36
rect 63 26 66 102
rect 75 96 80 102
rect 101 75 127 78
rect 49 23 66 26
rect 73 22 76 27
rect 84 17 89 36
rect 107 69 112 75
rect 14 14 89 17
rect 14 3 19 14
rect 38 5 41 10
rect 49 2 54 14
rect 84 13 89 14
rect 116 15 121 29
rect 73 5 76 10
rect 84 8 108 13
rect 116 10 127 15
rect 84 2 89 8
rect 116 2 121 10
rect 5 -42 10 -37
rect 40 -42 45 -38
rect 75 -42 80 -38
rect 107 -42 112 -38
rect 5 -45 112 -42
<< metal2 >>
rect 70 14 73 27
rect -1 11 73 14
rect 70 5 73 11
<< metal3 >>
rect 35 18 38 27
rect -1 15 38 18
rect 35 5 38 15
<< pad >>
rect 35 22 41 27
rect 70 22 76 27
rect 35 5 41 10
rect 70 5 76 10
<< labels >>
rlabel metal1 40 -45 45 -38 1 gnd!
rlabel metal1 101 75 127 78 1 vdd!
rlabel metal3 0 16 0 16 3 b
rlabel metal1 0 21 0 21 3 a
rlabel metal1 117 13 117 13 1 out
rlabel metal2 0 12 0 12 3 c
rlabel metal1 -1 102 25 105 5 vdd!
rlabel metal1 34 102 60 105 5 vdd!
rlabel metal1 69 102 95 105 5 vdd!
<< end >>
