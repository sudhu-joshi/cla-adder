magic
tech scmos
timestamp 1731965118
<< nwell >>
rect -58 219 -6 245
rect -58 187 -6 213
rect 74 212 126 238
rect -58 155 -6 181
rect 74 180 126 206
rect 78 145 130 171
rect -58 91 -6 117
rect -58 59 -6 85
rect 74 84 126 110
rect -58 27 -6 53
rect 74 52 126 78
rect 78 17 130 43
rect -58 -37 -6 -11
rect -58 -69 -6 -43
rect 74 -44 126 -18
rect -58 -101 -6 -75
rect 74 -76 126 -50
rect 78 -111 130 -85
rect -58 -165 -6 -139
rect -58 -197 -6 -171
rect 74 -172 126 -146
rect -58 -229 -6 -203
rect 74 -204 126 -178
rect 78 -239 130 -213
<< ntransistor >>
rect -120 231 -80 233
rect 13 224 53 226
rect -123 199 -83 201
rect 13 192 53 194
rect -119 167 -79 169
rect 13 157 53 159
rect -120 103 -80 105
rect 13 96 53 98
rect -123 71 -83 73
rect 13 64 53 66
rect -119 39 -79 41
rect 13 29 53 31
rect -120 -25 -80 -23
rect 13 -32 53 -30
rect -123 -57 -83 -55
rect 13 -64 53 -62
rect -119 -89 -79 -87
rect 13 -99 53 -97
rect -120 -153 -80 -151
rect 13 -160 53 -158
rect -123 -185 -83 -183
rect 13 -192 53 -190
rect -119 -217 -79 -215
rect 13 -227 53 -225
<< ptransistor >>
rect -52 231 -12 233
rect 80 224 120 226
rect -52 199 -12 201
rect 80 192 120 194
rect -52 167 -12 169
rect 84 157 124 159
rect -52 103 -12 105
rect 80 96 120 98
rect -52 71 -12 73
rect 80 64 120 66
rect -52 39 -12 41
rect 84 29 124 31
rect -52 -25 -12 -23
rect 80 -32 120 -30
rect -52 -57 -12 -55
rect 80 -64 120 -62
rect -52 -89 -12 -87
rect 84 -99 124 -97
rect -52 -153 -12 -151
rect 80 -160 120 -158
rect -52 -185 -12 -183
rect 80 -192 120 -190
rect -52 -217 -12 -215
rect 84 -227 124 -225
<< ndiffusion >>
rect -120 233 -80 234
rect -120 230 -80 231
rect 13 226 53 227
rect 13 223 53 224
rect -123 201 -83 202
rect -123 198 -83 199
rect 13 194 53 195
rect 13 191 53 192
rect -119 169 -79 170
rect -119 166 -79 167
rect 13 159 53 160
rect 13 156 53 157
rect -120 105 -80 106
rect -120 102 -80 103
rect 13 98 53 99
rect 13 95 53 96
rect -123 73 -83 74
rect -123 70 -83 71
rect 13 66 53 67
rect 13 63 53 64
rect -119 41 -79 42
rect -119 38 -79 39
rect 13 31 53 32
rect 13 28 53 29
rect -120 -23 -80 -22
rect -120 -26 -80 -25
rect 13 -30 53 -29
rect 13 -33 53 -32
rect -123 -55 -83 -54
rect -123 -58 -83 -57
rect 13 -62 53 -61
rect 13 -65 53 -64
rect -119 -87 -79 -86
rect -119 -90 -79 -89
rect 13 -97 53 -96
rect 13 -100 53 -99
rect -120 -151 -80 -150
rect -120 -154 -80 -153
rect 13 -158 53 -157
rect 13 -161 53 -160
rect -123 -183 -83 -182
rect -123 -186 -83 -185
rect 13 -190 53 -189
rect 13 -193 53 -192
rect -119 -215 -79 -214
rect -119 -218 -79 -217
rect 13 -225 53 -224
rect 13 -228 53 -227
<< pdiffusion >>
rect -52 233 -12 234
rect -52 230 -12 231
rect 80 226 120 227
rect 80 223 120 224
rect -52 201 -12 202
rect -52 198 -12 199
rect 80 194 120 195
rect 80 191 120 192
rect -52 169 -12 170
rect -52 166 -12 167
rect 84 159 124 160
rect 84 156 124 157
rect -52 105 -12 106
rect -52 102 -12 103
rect 80 98 120 99
rect 80 95 120 96
rect -52 73 -12 74
rect -52 70 -12 71
rect 80 66 120 67
rect 80 63 120 64
rect -52 41 -12 42
rect -52 38 -12 39
rect 84 31 124 32
rect 84 28 124 29
rect -52 -23 -12 -22
rect -52 -26 -12 -25
rect 80 -30 120 -29
rect 80 -33 120 -32
rect -52 -55 -12 -54
rect -52 -58 -12 -57
rect 80 -62 120 -61
rect 80 -65 120 -64
rect -52 -87 -12 -86
rect -52 -90 -12 -89
rect 84 -97 124 -96
rect 84 -100 124 -99
rect -52 -151 -12 -150
rect -52 -154 -12 -153
rect 80 -158 120 -157
rect 80 -161 120 -160
rect -52 -183 -12 -182
rect -52 -186 -12 -185
rect 80 -190 120 -189
rect 80 -193 120 -192
rect -52 -215 -12 -214
rect -52 -218 -12 -217
rect 84 -225 124 -224
rect 84 -228 124 -227
<< ndcontact >>
rect -120 234 -80 239
rect -120 225 -80 230
rect 13 227 53 232
rect 13 218 53 223
rect -123 202 -83 207
rect -123 193 -83 198
rect 13 195 53 200
rect 13 186 53 191
rect -119 170 -79 175
rect -119 161 -79 166
rect 13 160 53 165
rect 13 151 53 156
rect -120 106 -80 111
rect -120 97 -80 102
rect 13 99 53 104
rect 13 90 53 95
rect -123 74 -83 79
rect -123 65 -83 70
rect 13 67 53 72
rect 13 58 53 63
rect -119 42 -79 47
rect -119 33 -79 38
rect 13 32 53 37
rect 13 23 53 28
rect -120 -22 -80 -17
rect -120 -31 -80 -26
rect 13 -29 53 -24
rect 13 -38 53 -33
rect -123 -54 -83 -49
rect -123 -63 -83 -58
rect 13 -61 53 -56
rect 13 -70 53 -65
rect -119 -86 -79 -81
rect -119 -95 -79 -90
rect 13 -96 53 -91
rect 13 -105 53 -100
rect -120 -150 -80 -145
rect -120 -159 -80 -154
rect 13 -157 53 -152
rect 13 -166 53 -161
rect -123 -182 -83 -177
rect -123 -191 -83 -186
rect 13 -189 53 -184
rect 13 -198 53 -193
rect -119 -214 -79 -209
rect -119 -223 -79 -218
rect 13 -224 53 -219
rect 13 -233 53 -228
<< pdcontact >>
rect -52 234 -12 239
rect -52 225 -12 230
rect 80 227 120 232
rect 80 218 120 223
rect -52 202 -12 207
rect -52 193 -12 198
rect 80 195 120 200
rect 80 186 120 191
rect -52 170 -12 175
rect -52 161 -12 166
rect 84 160 124 165
rect 84 151 124 156
rect -52 106 -12 111
rect -52 97 -12 102
rect 80 99 120 104
rect 80 90 120 95
rect -52 74 -12 79
rect -52 65 -12 70
rect 80 67 120 72
rect 80 58 120 63
rect -52 42 -12 47
rect -52 33 -12 38
rect 84 32 124 37
rect 84 23 124 28
rect -52 -22 -12 -17
rect -52 -31 -12 -26
rect 80 -29 120 -24
rect 80 -38 120 -33
rect -52 -54 -12 -49
rect -52 -63 -12 -58
rect 80 -61 120 -56
rect 80 -70 120 -65
rect -52 -86 -12 -81
rect -52 -95 -12 -90
rect 84 -96 124 -91
rect 84 -105 124 -100
rect -52 -150 -12 -145
rect -52 -159 -12 -154
rect 80 -157 120 -152
rect 80 -166 120 -161
rect -52 -182 -12 -177
rect -52 -191 -12 -186
rect 80 -189 120 -184
rect 80 -198 120 -193
rect -52 -214 -12 -209
rect -52 -223 -12 -218
rect 84 -224 124 -219
rect 84 -233 124 -228
<< polysilicon >>
rect -123 231 -120 233
rect -80 231 -52 233
rect -12 231 -8 233
rect 10 224 13 226
rect 53 224 80 226
rect 120 224 124 226
rect -126 199 -123 201
rect -83 199 -74 201
rect -67 199 -52 201
rect -12 199 -8 201
rect 10 192 13 194
rect 53 192 80 194
rect 120 192 124 194
rect -122 167 -119 169
rect -79 167 -52 169
rect -12 167 -8 169
rect 10 157 13 159
rect 53 157 61 159
rect 68 157 84 159
rect 124 157 128 159
rect -123 103 -120 105
rect -80 103 -52 105
rect -12 103 -8 105
rect 10 96 13 98
rect 53 96 80 98
rect 120 96 124 98
rect -126 71 -123 73
rect -83 71 -74 73
rect -67 71 -52 73
rect -12 71 -8 73
rect 10 64 13 66
rect 53 64 80 66
rect 120 64 124 66
rect -122 39 -119 41
rect -79 39 -52 41
rect -12 39 -8 41
rect 10 29 13 31
rect 53 29 61 31
rect 68 29 84 31
rect 124 29 128 31
rect -123 -25 -120 -23
rect -80 -25 -52 -23
rect -12 -25 -8 -23
rect 10 -32 13 -30
rect 53 -32 80 -30
rect 120 -32 124 -30
rect -126 -57 -123 -55
rect -83 -57 -74 -55
rect -67 -57 -52 -55
rect -12 -57 -8 -55
rect 10 -64 13 -62
rect 53 -64 80 -62
rect 120 -64 124 -62
rect -122 -89 -119 -87
rect -79 -89 -52 -87
rect -12 -89 -8 -87
rect 10 -99 13 -97
rect 53 -99 61 -97
rect 68 -99 84 -97
rect 124 -99 128 -97
rect -123 -153 -120 -151
rect -80 -153 -52 -151
rect -12 -153 -8 -151
rect 10 -160 13 -158
rect 53 -160 80 -158
rect 120 -160 124 -158
rect -126 -185 -123 -183
rect -83 -185 -74 -183
rect -67 -185 -52 -183
rect -12 -185 -8 -183
rect 10 -192 13 -190
rect 53 -192 80 -190
rect 120 -192 124 -190
rect -122 -217 -119 -215
rect -79 -217 -52 -215
rect -12 -217 -8 -215
rect 10 -227 13 -225
rect 53 -227 61 -225
rect 68 -227 84 -225
rect 124 -227 128 -225
<< polycontact >>
rect -66 233 -61 238
rect 66 226 71 231
rect -80 201 -75 206
rect -66 201 -61 206
rect 57 194 62 199
rect -71 169 -66 174
rect 56 159 60 163
rect 71 159 76 164
rect -66 105 -61 110
rect 66 98 71 103
rect -80 73 -75 78
rect -66 73 -61 78
rect 57 66 62 71
rect -71 41 -66 46
rect 56 31 60 35
rect 71 31 76 36
rect -66 -23 -61 -18
rect 66 -30 71 -25
rect -80 -55 -75 -50
rect -66 -55 -61 -50
rect 57 -62 62 -57
rect -71 -87 -66 -82
rect 56 -97 60 -93
rect 71 -97 76 -92
rect -66 -151 -61 -146
rect 66 -158 71 -153
rect -80 -183 -75 -178
rect -66 -183 -61 -178
rect 57 -190 62 -185
rect -71 -215 -66 -210
rect 56 -225 60 -221
rect 71 -225 76 -220
<< metal1 >>
rect -134 234 -120 239
rect -66 238 -61 244
rect -6 239 0 245
rect -134 175 -130 234
rect -12 234 0 239
rect -80 222 -76 230
rect -127 218 -76 222
rect -66 225 -52 230
rect -66 219 -61 225
rect -127 202 -123 218
rect -72 214 -61 219
rect -80 206 -75 209
rect -72 198 -69 214
rect -66 206 -61 209
rect -6 207 0 234
rect 3 227 13 232
rect 66 231 71 237
rect 126 232 132 238
rect 3 218 7 227
rect 120 227 132 232
rect 53 218 80 223
rect 66 212 71 218
rect 126 212 132 227
rect -12 202 0 207
rect -83 193 -52 198
rect -134 170 -119 175
rect -71 174 -66 193
rect -6 175 0 202
rect 3 207 71 212
rect 3 200 6 207
rect 3 195 13 200
rect 57 199 62 202
rect 3 179 6 195
rect 120 195 131 200
rect 53 186 80 191
rect 3 175 60 179
rect -12 170 0 175
rect -79 161 -52 166
rect -71 139 -66 161
rect -6 155 0 170
rect 8 160 13 165
rect 56 163 60 175
rect 63 156 66 186
rect 71 164 76 167
rect 124 160 135 165
rect 53 151 84 156
rect 66 145 71 151
rect -134 106 -120 111
rect -66 110 -61 116
rect -6 111 0 117
rect -134 47 -130 106
rect -12 106 0 111
rect -80 94 -76 102
rect -127 90 -76 94
rect -66 97 -52 102
rect -66 91 -61 97
rect -127 74 -123 90
rect -72 86 -61 91
rect -80 78 -75 81
rect -72 70 -69 86
rect -66 78 -61 81
rect -6 79 0 106
rect 3 99 13 104
rect 66 103 71 109
rect 126 104 132 110
rect 3 90 7 99
rect 120 99 132 104
rect 53 90 80 95
rect 66 84 71 90
rect 126 84 132 99
rect -12 74 0 79
rect -83 65 -52 70
rect -134 42 -119 47
rect -71 46 -66 65
rect -6 47 0 74
rect 3 79 71 84
rect 3 72 6 79
rect 3 67 13 72
rect 57 71 62 74
rect 3 51 6 67
rect 120 67 131 72
rect 53 58 80 63
rect 3 47 60 51
rect -12 42 0 47
rect -79 33 -52 38
rect -71 11 -66 33
rect -6 27 0 42
rect 8 32 13 37
rect 56 35 60 47
rect 63 28 66 58
rect 71 36 76 39
rect 124 32 135 37
rect 53 23 84 28
rect 66 17 71 23
rect -134 -22 -120 -17
rect -66 -18 -61 -12
rect -6 -17 0 -11
rect -134 -81 -130 -22
rect -12 -22 0 -17
rect -80 -34 -76 -26
rect -127 -38 -76 -34
rect -66 -31 -52 -26
rect -66 -37 -61 -31
rect -127 -54 -123 -38
rect -72 -42 -61 -37
rect -80 -50 -75 -47
rect -72 -58 -69 -42
rect -66 -50 -61 -47
rect -6 -49 0 -22
rect 3 -29 13 -24
rect 66 -25 71 -19
rect 126 -24 132 -18
rect 3 -38 7 -29
rect 120 -29 132 -24
rect 53 -38 80 -33
rect 66 -44 71 -38
rect 126 -44 132 -29
rect -12 -54 0 -49
rect -83 -63 -52 -58
rect -134 -86 -119 -81
rect -71 -82 -66 -63
rect -6 -81 0 -54
rect 3 -49 71 -44
rect 3 -56 6 -49
rect 3 -61 13 -56
rect 57 -57 62 -54
rect 3 -77 6 -61
rect 120 -61 131 -56
rect 53 -70 80 -65
rect 3 -81 60 -77
rect -12 -86 0 -81
rect -79 -95 -52 -90
rect -71 -117 -66 -95
rect -6 -101 0 -86
rect 8 -96 13 -91
rect 56 -93 60 -81
rect 63 -100 66 -70
rect 71 -92 76 -89
rect 124 -96 135 -91
rect 53 -105 84 -100
rect 66 -111 71 -105
rect -134 -150 -120 -145
rect -66 -146 -61 -140
rect -6 -145 0 -139
rect -134 -209 -130 -150
rect -12 -150 0 -145
rect -80 -162 -76 -154
rect -127 -166 -76 -162
rect -66 -159 -52 -154
rect -66 -165 -61 -159
rect -127 -182 -123 -166
rect -72 -170 -61 -165
rect -80 -178 -75 -175
rect -72 -186 -69 -170
rect -66 -178 -61 -175
rect -6 -177 0 -150
rect 3 -157 13 -152
rect 66 -153 71 -147
rect 126 -152 132 -146
rect 3 -166 7 -157
rect 120 -157 132 -152
rect 53 -166 80 -161
rect 66 -172 71 -166
rect 126 -172 132 -157
rect -12 -182 0 -177
rect -83 -191 -52 -186
rect -134 -214 -119 -209
rect -71 -210 -66 -191
rect -6 -209 0 -182
rect 3 -177 71 -172
rect 3 -184 6 -177
rect 3 -189 13 -184
rect 57 -185 62 -182
rect 3 -205 6 -189
rect 120 -189 131 -184
rect 53 -198 80 -193
rect 3 -209 60 -205
rect -12 -214 0 -209
rect -79 -223 -52 -218
rect -71 -245 -66 -223
rect -6 -229 0 -214
rect 8 -224 13 -219
rect 56 -221 60 -209
rect 63 -228 66 -198
rect 71 -220 76 -217
rect 124 -224 135 -219
rect 53 -233 84 -228
rect 66 -239 71 -233
rect -138 -273 -114 -266
<< metal2 >>
rect -134 250 71 253
rect -66 241 -61 250
rect 66 245 71 250
rect 66 241 138 245
rect 66 234 71 241
rect 134 200 138 241
rect 131 195 138 200
rect 134 179 138 195
rect 71 176 138 179
rect 71 167 76 176
rect -134 122 71 125
rect -66 113 -61 122
rect 66 117 71 122
rect 66 113 138 117
rect 66 106 71 113
rect 134 72 138 113
rect 131 67 138 72
rect 134 51 138 67
rect 71 48 138 51
rect 71 39 76 48
rect -134 -6 71 -3
rect -66 -15 -61 -6
rect 66 -11 71 -6
rect 66 -15 138 -11
rect 66 -22 71 -15
rect 134 -56 138 -15
rect 131 -61 138 -56
rect 134 -77 138 -61
rect 71 -80 138 -77
rect 71 -89 76 -80
rect -134 -134 71 -131
rect -66 -143 -61 -134
rect 66 -139 71 -134
rect 66 -143 138 -139
rect 66 -150 71 -143
rect 134 -184 138 -143
rect 131 -189 138 -184
rect 134 -205 138 -189
rect 71 -208 138 -205
rect 71 -217 76 -208
<< metal3 >>
rect -134 246 62 249
rect -74 212 -69 246
rect -80 209 -61 212
rect 57 211 62 246
rect 57 207 143 211
rect 57 202 62 207
rect 140 175 143 207
rect 60 172 143 175
rect 1 169 63 172
rect 1 165 5 169
rect 140 165 143 172
rect 1 160 8 165
rect 135 160 143 165
rect -134 118 62 121
rect -74 84 -69 118
rect -80 81 -61 84
rect 57 83 62 118
rect 57 79 143 83
rect 57 74 62 79
rect 140 47 143 79
rect 60 44 143 47
rect 1 41 63 44
rect 1 37 5 41
rect 140 37 143 44
rect 1 32 8 37
rect 135 32 143 37
rect -134 -10 62 -7
rect -74 -44 -69 -10
rect -80 -47 -61 -44
rect 57 -45 62 -10
rect 57 -49 143 -45
rect 57 -54 62 -49
rect 140 -81 143 -49
rect 60 -84 143 -81
rect 1 -87 63 -84
rect 1 -91 5 -87
rect 140 -91 143 -84
rect 1 -96 8 -91
rect 135 -96 143 -91
rect -134 -138 62 -135
rect -74 -172 -69 -138
rect -80 -175 -61 -172
rect 57 -173 62 -138
rect 57 -177 143 -173
rect 57 -182 62 -177
rect 140 -209 143 -177
rect 60 -212 143 -209
rect 1 -215 63 -212
rect 1 -219 5 -215
rect 140 -219 143 -212
rect 1 -224 8 -219
rect 135 -224 143 -219
<< metal5 >>
rect 66 142 71 145
rect 66 137 143 142
rect 66 14 71 17
rect 66 9 143 14
rect 66 -114 71 -111
rect 66 -119 143 -114
rect 66 -242 71 -239
rect 66 -247 143 -242
<< metal6 >>
rect -71 131 143 136
rect -71 3 143 8
rect -71 -125 143 -120
rect -71 -253 143 -248
<< pad >>
rect -66 238 -61 244
rect 66 231 71 237
rect -80 206 -75 212
rect -66 206 -61 212
rect 57 199 62 204
rect 128 195 134 200
rect 5 160 11 165
rect 71 164 76 170
rect 132 160 138 165
rect 66 142 71 148
rect -71 136 -66 142
rect -66 110 -61 116
rect 66 103 71 109
rect -80 78 -75 84
rect -66 78 -61 84
rect 57 71 62 76
rect 128 67 134 72
rect 5 32 11 37
rect 71 36 76 42
rect 132 32 138 37
rect 66 14 71 20
rect -71 8 -66 14
rect -66 -18 -61 -12
rect 66 -25 71 -19
rect -80 -50 -75 -44
rect -66 -50 -61 -44
rect 57 -57 62 -52
rect 128 -61 134 -56
rect 5 -96 11 -91
rect 71 -92 76 -86
rect 132 -96 138 -91
rect 66 -114 71 -108
rect -71 -120 -66 -114
rect -66 -146 -61 -140
rect 66 -153 71 -147
rect -80 -178 -75 -172
rect -66 -178 -61 -172
rect 57 -185 62 -180
rect 128 -189 134 -184
rect 5 -224 11 -219
rect 71 -220 76 -214
rect 132 -224 138 -219
rect 66 -242 71 -236
rect -71 -248 -66 -242
<< labels >>
rlabel metal1 126 84 132 110 1 vdd!
rlabel metal1 3 90 7 104 1 gnd!
rlabel metal1 -134 42 -130 111 3 gnd!
rlabel metal1 -6 27 0 117 1 vdd!
rlabel metal1 126 212 132 238 1 vdd!
rlabel metal1 3 218 7 232 1 gnd!
rlabel metal1 -134 170 -130 239 3 gnd!
rlabel metal1 -6 155 0 245 1 vdd!
rlabel metal1 -6 -101 0 -11 1 vdd!
rlabel metal1 -134 -86 -130 -17 3 gnd!
rlabel metal1 3 -38 7 -24 1 gnd!
rlabel metal1 126 -44 132 -18 1 vdd!
rlabel metal1 -6 -229 0 -139 1 vdd!
rlabel metal1 -134 -214 -130 -145 3 gnd!
rlabel metal1 3 -166 7 -152 1 gnd!
rlabel metal1 126 -172 132 -146 1 vdd!
rlabel metal6 -71 -253 143 -248 1 g0
rlabel metal5 66 -247 143 -242 1 p0
rlabel metal6 -71 -125 143 -120 1 g1
rlabel metal5 66 -119 143 -114 1 p1
rlabel metal3 57 -54 62 -7 1 b1
rlabel metal2 -134 -6 71 -3 1 a1
rlabel metal3 -134 -138 62 -135 1 b0
rlabel metal2 -134 -134 71 -131 1 a0
rlabel metal3 -134 -10 62 -7 1 b1
rlabel metal3 -134 118 62 121 1 b2
rlabel metal2 -134 122 71 125 1 a2
rlabel metal6 -71 3 143 8 1 g2
rlabel metal5 66 9 143 14 1 p2
rlabel metal6 -71 131 143 136 1 g3
rlabel metal5 66 137 143 142 1 p3
rlabel metal2 -134 250 71 253 5 a3
rlabel metal3 -134 246 62 249 1 b3
rlabel metal1 -138 -273 -114 -266 1 c0
<< end >>
