* SPICE3 file created from final_cla.ext - technology: scmos

.option scale=0.09u

M1000 a_148_74# g0 vdd w_166_68# pfet w=40 l=2
+  ad=720 pd=276 as=17634 ps=6694
M1001 vdd a1 a_n266_n63# w_n201_n37# pfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1002 a_44_n176# p1 gnd Gnd nfet w=60 l=2
+  ad=720 pd=264 as=14160 ps=5368
M1003 a_148_n14# p2 gnd Gnd nfet w=60 l=2
+  ad=720 pd=264 as=0 ps=0
M1004 a_279_n316# a_240_n171# gnd Gnd nfet w=40 l=2
+  ad=720 pd=276 as=0 ps=0
M1005 c2 a_279_n316# gnd Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1006 a_676_n97# p2 gnd Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1007 a_507_198# a_426_70# a_472_198# w_493_192# pfet w=199 l=2
+  ad=2388 pd=820 as=2388 ps=820
M1008 c3 a_441_n306# gnd Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1009 a_418_n118# a_290_n49# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1010 a_244_7# a_148_74# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1011 a_290_n49# p2 vdd w_372_n55# pfet w=40 l=2
+  ad=960 pd=368 as=0 ps=0
M1012 a_n266_n183# b0 a_n266_n191# Gnd nfet w=40 l=2
+  ad=480 pd=184 as=240 ps=92
M1013 a_322_n165# c0 a_290_n159# Gnd nfet w=80 l=2
+  ad=960 pd=344 as=960 ps=344
M1014 vdd a1 a_n133_n99# w_n69_n44# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1015 a_140_n155# a_44_n88# vdd w_126_n94# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1016 a_542_198# a_241_164# a_507_198# w_528_192# pfet w=199 l=2
+  ad=2388 pd=820 as=0 ps=0
M1017 a_44_n241# p0 vdd w_30_n247# pfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1018 a_34_206# p3 vdd w_20_200# pfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1019 a_298_139# p2 vdd w_380_133# pfet w=40 l=2
+  ad=960 pd=368 as=0 ps=0
M1020 c3 a_441_n306# vdd w_564_n242# pfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1021 b0 a_n133_n227# p0 Gnd nfet w=40 l=2
+  ad=240 pd=92 as=480 ps=184
M1022 b3 a_n133_157# p3 Gnd nfet w=40 l=2
+  ad=240 pd=92 as=480 ps=184
M1023 vdd a2 a_n133_29# w_n69_84# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1024 a_n133_29# b2 p2 Gnd nfet w=40 l=2
+  ad=480 pd=184 as=480 ps=184
M1025 a_298_29# p3 gnd Gnd nfet w=80 l=2
+  ad=960 pd=344 as=0 ps=0
M1026 vdd b3 a_n266_193# w_n201_187# pfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1027 a_472_117# a_605_159# gnd Gnd nfet w=40 l=2
+  ad=1200 pd=460 as=0 ps=0
M1028 a_n266_n55# b1 a_n266_n63# Gnd nfet w=40 l=2
+  ad=480 pd=184 as=240 ps=92
M1029 a_44_n309# p0 gnd Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1030 s0 c0 p0 w_671_n328# pfet w=40 l=2
+  ad=480 pd=184 as=720 ps=276
M1031 s1 c1 p1 w_671_n183# pfet w=40 l=2
+  ad=480 pd=184 as=720 ps=276
M1032 a_145_231# p2 vdd w_195_225# pfet w=40 l=2
+  ad=720 pd=276 as=0 ps=0
M1033 a_426_70# a_298_139# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1034 a_n133_n99# b1 p1 Gnd nfet w=40 l=2
+  ad=480 pd=184 as=480 ps=184
M1035 a_476_n229# a_244_7# a_441_n229# w_462_n235# pfet w=80 l=2
+  ad=960 pd=344 as=960 ps=344
M1036 a_44_n88# p1 vdd w_30_n94# pfet w=40 l=2
+  ad=720 pd=276 as=0 ps=0
M1037 b3 a3 p3 w_n65_145# pfet w=40 l=2
+  ad=240 pd=92 as=720 ps=276
M1038 a_106_n9# a_42_58# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1039 a_44_n88# p0 a_76_n182# Gnd nfet w=60 l=2
+  ad=360 pd=132 as=720 ps=264
M1040 a_459_n85# p3 gnd Gnd nfet w=100 l=2
+  ad=1200 pd=424 as=0 ps=0
M1041 gnd a2 a_n266_73# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1042 a_145_231# p3 vdd w_131_225# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 s2 c2 p2 w_694_n36# pfet w=40 l=2
+  ad=480 pd=184 as=720 ps=276
M1044 a_290_n49# p0 vdd w_276_n55# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 vdd a3 a_n133_157# w_n69_212# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1046 a_98_139# a_34_206# vdd w_84_200# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1047 a_241_164# a_145_231# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1048 s1 c1 a_653_n244# Gnd nfet w=40 l=2
+  ad=480 pd=184 as=480 ps=184
M1049 gnd a0 a_n133_n227# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1050 a_472_117# a_98_139# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 a_676_48# p3 vdd w_662_109# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1052 a_511_n229# a_106_n9# a_476_n229# w_497_n235# pfet w=80 l=2
+  ad=960 pd=344 as=0 ps=0
M1053 a_298_139# p3 vdd w_284_133# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 a_42_58# g1 a_42_n10# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=480 ps=184
M1055 a_279_n316# a_140_n155# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 c4 a_472_117# vdd w_630_183# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1057 a_148_74# p1 a_180_n20# Gnd nfet w=60 l=2
+  ad=360 pd=132 as=720 ps=264
M1058 a_459_51# p1 vdd w_509_45# pfet w=40 l=2
+  ad=1200 pd=460 as=0 ps=0
M1059 a_279_n316# a_140_n155# a_314_n243# w_335_n249# pfet w=60 l=2
+  ad=360 pd=132 as=720 ps=264
M1060 s2 c2 a_676_n97# Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1061 a_240_n171# a_176_n104# vdd w_226_n110# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1062 a_441_n306# a_418_n118# gnd Gnd nfet w=40 l=2
+  ad=960 pd=368 as=0 ps=0
M1063 a_523_n91# p1 a_491_n91# Gnd nfet w=100 l=2
+  ad=1200 pd=424 as=1200 ps=424
M1064 a_177_137# g1 a_145_143# Gnd nfet w=60 l=2
+  ad=720 pd=264 as=720 ps=264
M1065 a_42_58# p2 vdd w_28_52# pfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1066 a_290_n159# p0 gnd Gnd nfet w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 a_244_7# a_148_74# vdd w_230_68# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1068 a_362_23# p1 a_330_23# Gnd nfet w=80 l=2
+  ad=960 pd=344 as=960 ps=344
M1069 a_148_74# p2 vdd w_134_68# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 vdd b0 a_n266_n191# w_n201_n197# pfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1071 a_418_n118# a_290_n49# vdd w_404_n55# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1072 a_140_n320# g0 a_140_n252# w_163_n258# pfet w=40 l=2
+  ad=240 pd=92 as=480 ps=184
M1073 a_290_n49# p2 a_354_n165# Gnd nfet w=80 l=2
+  ad=480 pd=172 as=960 ps=344
M1074 a_472_117# a_426_70# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 c1 a_140_n320# vdd w_195_n258# pfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1076 a_108_n308# a_44_n241# vdd w_94_n247# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1077 vdd a3 a_n266_193# w_n201_219# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 a_n133_157# b3 p3 Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1079 gnd a_n266_193# g3 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1080 s1 a_653_n244# c1 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1081 s2 a_676_n97# c2 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 a_240_n171# a_176_n104# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1083 a_176_n172# p1 gnd Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1084 a_34_206# g2 a_34_138# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=480 ps=184
M1085 a_472_198# g3 vdd w_458_192# pfet w=199 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 a_106_n9# a_42_58# vdd w_92_52# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1087 vdd b1 a_n266_n63# w_n201_n69# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 a_290_n49# p1 vdd w_340_n55# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 a_426_70# a_298_139# vdd w_412_133# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1090 a_140_n320# g0 gnd Gnd nfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1091 gnd a1 a_n266_n55# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 a_140_n252# a_108_n308# vdd w_126_n258# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 vdd a0 a_n133_n227# w_n69_n172# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1094 a_44_n88# p0 vdd w_94_n94# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 gnd a0 a_n266_n183# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 a_472_117# a_241_164# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 a_441_n306# g2 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1098 s3 p3 c3 w_729_113# pfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1099 s0 c0 a_653_n389# Gnd nfet w=40 l=2
+  ad=480 pd=184 as=480 ps=184
M1100 a_653_n389# p0 vdd w_639_n328# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1101 a_653_n244# p1 vdd w_639_n183# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1102 vdd a_n266_65# g2 w_n201_27# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1103 s1 p1 c1 w_706_n179# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 a_298_139# p1 vdd w_348_133# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 a_459_51# p0 vdd w_573_45# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 a1 b1 p1 w_n69_n76# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1107 a_n133_n227# b0 p0 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 a_176_n104# g0 a_176_n172# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1109 a_472_117# g3 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 a_140_n320# a_108_n308# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 a_459_51# p0 a_555_n91# Gnd nfet w=100 l=2
+  ad=600 pd=212 as=1200 ps=424
M1112 a_459_51# c0 vdd w_477_45# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 a_279_n316# g1 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 a_314_n243# g1 a_279_n243# w_300_n249# pfet w=60 l=2
+  ad=0 pd=0 as=720 ps=264
M1115 s2 p2 c2 w_729_n32# pfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1116 a_76_n182# c0 a_44_n176# Gnd nfet w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 gnd a2 a_n133_29# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 a_605_159# a_459_51# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1119 s0 a_653_n389# c0 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1120 a_653_n244# p1 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 s3 c3 a_676_48# Gnd nfet w=40 l=2
+  ad=480 pd=184 as=480 ps=184
M1122 gnd a_n266_n63# g1 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1123 s3 c3 p3 w_694_109# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 a_176_n104# p1 vdd w_162_n110# pfet w=40 l=2
+  ad=480 pd=184 as=0 ps=0
M1125 a2 b2 p2 w_n69_52# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1126 a_44_n241# c0 a_44_n309# Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1127 a_176_n104# g0 vdd w_194_n110# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 a_298_139# g0 vdd w_316_133# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 a_441_n229# g2 vdd w_427_n235# pfet w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 vdd a_n266_193# g3 w_n201_155# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1131 a_145_143# p3 gnd Gnd nfet w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 b2 a2 p2 w_n65_17# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1133 a0 b0 p0 w_n69_n204# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1134 a_34_206# g2 vdd w_52_200# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 a_145_231# p2 a_177_137# Gnd nfet w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1136 a_n266_73# b2 a_n266_65# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1137 a_279_n243# a_240_n171# vdd w_265_n249# pfet w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 a_441_n306# a_244_7# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 s3 a_676_48# c3 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 a_354_n165# p1 a_322_n165# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 a_605_159# a_459_51# vdd w_607_45# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1142 gnd a1 a_n133_n99# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 b1 a_n133_n99# p1 Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1144 vdd b2 a_n266_65# w_n201_59# pfet w=40 l=2
+  ad=0 pd=0 as=480 ps=184
M1145 c4 a_472_117# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1146 b0 a0 p0 w_n65_n239# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1147 a_472_117# a_605_159# a_577_198# w_598_192# pfet w=199 l=2
+  ad=1194 pd=410 as=2388 ps=820
M1148 a_180_n20# g0 a_148_n14# Gnd nfet w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1149 gnd a_n266_n191# g0 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1150 a_491_n91# c0 a_459_n85# Gnd nfet w=100 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 vdd a2 a_n266_65# w_n201_91# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 a3 b3 p3 w_n69_180# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1153 gnd a_n266_65# g2 Gnd nfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1154 s0 p0 c0 w_706_n324# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1155 a_44_n241# c0 vdd w_62_n247# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1156 c1 a_140_n320# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 a_241_164# a_145_231# vdd w_227_225# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1158 a_148_74# p1 vdd w_198_68# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 a_108_n308# a_44_n241# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1160 a_676_48# p3 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 a_98_139# a_34_206# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1162 a_44_n88# c0 vdd w_62_n94# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1163 b2 a_n133_29# p2 Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1164 a_330_23# g0 a_298_29# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 a_653_n389# p0 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 a_441_n306# a_106_n9# gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 b1 a1 p1 w_n65_n111# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1168 a_441_n306# a_418_n118# a_511_n229# w_532_n235# pfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1169 a_145_231# g1 vdd w_163_225# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 a_42_n10# p2 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 a_n266_201# b3 a_n266_193# Gnd nfet w=40 l=2
+  ad=480 pd=184 as=240 ps=92
M1172 a_290_n49# c0 vdd w_308_n55# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 c2 a_279_n316# vdd w_367_n256# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 gnd a3 a_n266_201# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 vdd a_n266_n191# g0 w_n201_n229# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1176 a_140_n155# a_44_n88# gnd Gnd nfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1177 vdd a_n266_n63# g1 w_n201_n101# pfet w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1178 a_577_198# a_98_139# a_542_198# w_563_192# pfet w=199 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 a_676_n97# p2 vdd w_662_n36# pfet w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1180 vdd a0 a_n266_n191# w_n201_n165# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 a_34_138# p3 gnd Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 gnd a3 a_n133_157# Gnd nfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 a_459_51# p2 vdd w_541_45# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 a_555_n91# p2 a_523_n91# Gnd nfet w=100 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 a_459_51# p3 vdd w_445_45# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 a_42_58# g1 vdd w_60_52# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 a_298_139# p2 a_362_23# Gnd nfet w=80 l=2
+  ad=480 pd=172 as=0 ps=0
C0 w_n201_59# a_n266_65# 0.07fF
C1 w_134_68# g0 0.01fF
C2 w_30_n94# vdd 0.09fF
C3 p1 a_298_139# 0.73fF
C4 w_230_68# a_148_74# 0.07fF
C5 w_92_52# a_42_58# 0.07fF
C6 w_372_n55# vdd 0.09fF
C7 g1 a_n266_n63# 0.07fF
C8 p1 a_180_n20# 0.08fF
C9 w_226_n110# vdd 0.09fF
C10 g0 a_298_29# 0.10fF
C11 a_n266_65# b2 0.48fF
C12 a_n266_n191# vdd 0.89fF
C13 g0 p0 0.18fF
C14 p1 c0 0.34fF
C15 a_298_139# a_362_23# 0.82fF
C16 w_694_n36# p2 0.07fF
C17 p1 a_44_n88# 0.07fF
C18 w_573_45# p0 0.07fF
C19 w_541_45# a_459_51# 0.07fF
C20 w_n65_n111# p1 0.07fF
C21 a_298_29# a_330_23# 0.82fF
C22 c3 s3 0.95fF
C23 a_491_n91# a_523_n91# 1.03fF
C24 w_n201_n37# a_n266_n63# 0.07fF
C25 w_340_n55# p1 0.07fF
C26 a_244_7# a_418_n118# 0.06fF
C27 c2 s2 0.95fF
C28 a_290_n159# a_279_n243# 0.15fF
C29 w_n65_n111# a1 0.07fF
C30 g0 a_n266_n191# 0.07fF
C31 a_76_n182# vdd 0.25fF
C32 a_44_n176# gnd 0.72fF
C33 c1 a_140_n320# 0.07fF
C34 a_44_n241# a_108_n308# 0.07fF
C35 p0 a0 0.55fF
C36 a_n266_n63# b1 0.48fF
C37 a_290_n49# a_418_n118# 0.07fF
C38 w_126_n258# a_108_n308# 0.07fF
C39 w_195_n258# c1 0.07fF
C40 w_308_n55# c0 0.07fF
C41 w_276_n55# p0 0.07fF
C42 w_265_n249# a_279_n243# 0.09fF
C43 a_108_n308# vdd 0.45fF
C44 w_162_n110# c0 0.01fF
C45 w_126_n94# a_140_n155# 0.07fF
C46 w_427_n235# a_441_n229# 0.11fF
C47 a_441_n229# vdd 0.90fF
C48 a_279_n243# gnd 0.02fF
C49 p2 a_676_n97# 0.08fF
C50 vdd a_653_n389# 0.45fF
C51 a_653_n244# gnd 0.47fF
C52 a0 a_n266_n191# 0.07fF
C53 w_639_n328# vdd 0.09fF
C54 g1 a_279_n243# 0.02fF
C55 w_163_225# vdd 0.09fF
C56 p1 a_491_n91# 0.10fF
C57 a_605_159# vdd 2.92fF
C58 a_426_70# gnd 0.51fF
C59 g0 a_108_n308# 0.04fF
C60 a_145_231# gnd 0.03fF
C61 w_n201_155# vdd 0.07fF
C62 w_458_192# g3 0.07fF
C63 w_630_183# vdd 0.09fF
C64 w_163_n258# g0 0.07fF
C65 c0 a_240_n171# 0.04fF
C66 a_98_139# a_605_159# 0.06fF
C67 a_241_164# p3 0.08fF
C68 w_227_225# a_145_231# 0.07fF
C69 w_60_52# vdd 0.09fF
C70 g1 a_145_231# 0.37fF
C71 p1 vdd 0.05fF
C72 c0 a_459_n85# 0.10fF
C73 a_290_n49# a_290_n159# 0.08fF
C74 p3 g2 0.00fF
C75 a_426_70# a_507_198# 0.05fF
C76 a_n266_n183# b0 0.07fF
C77 a_42_58# vdd 0.89fF
C78 a_176_n104# a_176_n172# 0.42fF
C79 c0 c1 0.66fF
C80 a_106_n9# a_441_n306# 0.83fF
C81 w_n69_212# a3 0.07fF
C82 w_n201_219# a_n266_193# 0.07fF
C83 w_607_45# vdd 0.09fF
C84 w_493_192# a_507_198# 0.23fF
C85 a_n266_193# b3 0.48fF
C86 c3 a_441_n306# 0.07fF
C87 a_244_7# gnd 0.51fF
C88 a_676_48# gnd 0.47fF
C89 p2 a_148_74# 0.07fF
C90 a_145_143# a_177_137# 0.62fF
C91 w_380_133# a_298_139# 0.07fF
C92 a_418_n118# a_511_n229# 0.04fF
C93 p2 a_106_n9# 0.07fF
C94 a_n133_n99# vdd 0.96fF
C95 a_472_198# a_472_117# 0.12fF
C96 p3 s3 0.55fF
C97 g0 p1 0.68fF
C98 a_418_n118# gnd 0.77fF
C99 p2 c3 0.60fF
C100 w_532_n235# a_418_n118# 0.07fF
C101 a_241_164# c0 0.08fF
C102 w_28_52# a_42_58# 0.07fF
C103 w_166_68# a_148_74# 0.07fF
C104 g2 c0 0.08fF
C105 w_308_n55# vdd 0.09fF
C106 p2 a_459_51# 0.20fF
C107 a2 b2 0.23fF
C108 w_162_n110# vdd 0.09fF
C109 a_148_74# a_106_n9# 0.03fF
C110 p1 a_330_23# 0.10fF
C111 a_44_n176# a_76_n182# 0.62fF
C112 w_729_113# s3 0.07fF
C113 w_477_45# a_459_51# 0.07fF
C114 a_244_7# p0 0.07fF
C115 a_n133_n227# gnd 0.47fF
C116 a_459_n85# a_491_n91# 1.03fF
C117 a_330_23# a_362_23# 0.82fF
C118 a1 a_n266_n63# 0.07fF
C119 p0 a_290_n49# 0.07fF
C120 w_n69_n172# vdd 0.09fF
C121 a_240_n171# vdd 0.45fF
C122 c0 a_176_n104# 0.08fF
C123 a_290_n159# gnd 0.93fF
C124 w_94_n247# a_44_n241# 0.07fF
C125 a_140_n320# a_140_n252# 0.45fF
C126 w_126_n94# c0 0.01fF
C127 w_94_n94# p0 0.07fF
C128 c1 vdd 0.45fF
C129 a_314_n243# a_279_n316# 0.77fF
C130 c2 gnd 0.41fF
C131 w_126_n94# a_44_n88# 0.07fF
C132 w_372_n55# a_290_n49# 0.07fF
C133 a_476_n229# a_441_n306# 0.12fF
C134 a_44_n309# gnd 0.69fF
C135 w_367_n256# a_279_n316# 0.07fF
C136 w_94_n247# vdd 0.09fF
C137 p2 a_555_n91# 0.01fF
C138 w_367_n256# vdd 0.09fF
C139 w_532_n235# a_511_n229# 0.13fF
C140 w_194_n110# a_176_n104# 0.07fF
C141 p0 a_n133_n227# 1.05fF
C142 a_241_164# vdd 0.45fF
C143 p1 a_354_n165# 0.01fF
C144 g2 vdd 0.41fF
C145 g1 gnd 0.48fF
C146 w_427_n235# g2 0.07fF
C147 w_n201_187# vdd 0.09fF
C148 w_380_133# vdd 0.09fF
C149 a_426_70# a_605_159# 0.21fF
C150 g3 p3 0.75fF
C151 a_241_164# a_98_139# 0.71fF
C152 a_n266_193# gnd 0.03fF
C153 w_195_225# p2 0.07fF
C154 w_163_225# a_145_231# 0.07fF
C155 c0 a_322_n165# 0.01fF
C156 p3 p2 0.05fF
C157 p1 a_653_n244# 0.08fF
C158 w_n69_n172# a0 0.07fF
C159 w_230_68# vdd 0.09fF
C160 a_106_n9# a_476_n229# 0.02fF
C161 a_244_7# a_441_n229# 0.02fF
C162 g3 a_472_198# 0.01fF
C163 g2 a_34_206# 0.48fF
C164 p1 m5_167_n48# 0.00fF
C165 a_459_51# a_555_n91# 1.03fF
C166 w_671_n183# p1 0.07fF
C167 c4 gnd 0.41fF
C168 p3 a_n133_157# 1.05fF
C169 w_n201_219# a3 0.07fF
C170 w_458_192# a_472_198# 0.23fF
C171 w_541_45# vdd 0.09fF
C172 w_n65_n239# p0 0.07fF
C173 w_497_n235# a_106_n9# 0.07fF
C174 a3 b3 0.23fF
C175 a_605_159# a_577_198# 0.02fF
C176 a_34_206# a_34_138# 0.42fF
C177 w_462_n235# a_244_7# 0.07fF
C178 a_98_139# a_472_117# 0.19fF
C179 a_145_231# a_177_137# 0.62fF
C180 w_598_192# a_577_198# 0.25fF
C181 w_n201_n101# vdd 0.09fF
C182 p2 a_298_139# 0.27fF
C183 g2 g0 0.04fF
C184 a_298_29# gnd 0.93fF
C185 w_316_133# a_298_139# 0.07fF
C186 w_348_133# p1 0.07fF
C187 g2 a_n266_65# 0.07fF
C188 p2 a_n133_29# 1.05fF
C189 w_n65_17# p2 0.07fF
C190 p3 c3 0.15fF
C191 w_706_n324# p0 0.07fF
C192 a_176_n104# vdd 0.89fF
C193 w_198_68# p1 0.07fF
C194 w_n201_59# b2 0.07fF
C195 w_n69_84# a_n133_29# 0.07fF
C196 w_126_n94# vdd 0.09fF
C197 g1 p0 0.18fF
C198 p3 a_459_51# 0.07fF
C199 p2 c0 0.26fF
C200 w_n201_n197# b0 0.07fF
C201 w_509_45# p1 0.07fF
C202 w_92_52# a_106_n9# 0.07fF
C203 a_n266_73# a_n266_65# 0.42fF
C204 p1 a_244_7# 0.13fF
C205 a_148_74# a_180_n20# 0.62fF
C206 a_n266_n191# gnd 0.03fF
C207 w_729_113# c3 0.07fF
C208 p1 a_290_n49# 0.73fF
C209 a_106_n9# a_180_n20# 0.25fF
C210 w_n69_n44# a1 0.07fF
C211 w_477_45# c0 0.07fF
C212 g0 a_176_n104# 0.48fF
C213 w_n201_n197# vdd 0.09fF
C214 w_126_n94# g0 0.19fF
C215 a_240_n171# a_279_n243# 0.01fF
C216 w_n69_n44# a_n133_n99# 0.07fF
C217 w_n201_n101# a_n266_n63# 0.07fF
C218 c0 a_459_51# 0.32fF
C219 c0 a_140_n155# 0.05fF
C220 a_n266_n55# a_n266_n63# 0.42fF
C221 w_30_n247# a_44_n241# 0.07fF
C222 w_62_n94# c0 0.08fF
C223 a_44_n88# a_140_n155# 0.07fF
C224 c1 a_653_n244# 0.40fF
C225 w_195_n258# a_140_n320# 0.07fF
C226 a_279_n243# a_314_n243# 0.69fF
C227 a_676_n97# vdd 0.45fF
C228 a_523_n91# gnd 0.25fF
C229 w_126_n258# a_140_n252# 0.07fF
C230 w_62_n94# a_44_n88# 0.07fF
C231 w_308_n55# a_290_n49# 0.07fF
C232 w_671_n183# c1 0.07fF
C233 w_30_n247# vdd 0.09fF
C234 w_335_n249# a_314_n243# 0.11fF
C235 a_140_n252# vdd 0.98fF
C236 a_108_n308# gnd 0.41fF
C237 w_226_n110# p0 0.02fF
C238 a_653_n244# s1 1.05fF
C239 w_497_n235# a_476_n229# 0.13fF
C240 w_639_n183# vdd 0.09fF
C241 vdd m1_163_n48# 0.03fF
C242 w_671_n183# s1 0.07fF
C243 w_564_n242# a_441_n306# 0.07fF
C244 a_653_n389# gnd 0.47fF
C245 g3 vdd 0.41fF
C246 w_671_n328# s0 0.07fF
C247 w_458_192# vdd 0.25fF
C248 a_605_159# gnd 2.91fF
C249 w_316_133# vdd 0.09fF
C250 a_n133_157# vdd 0.96fF
C251 a_426_70# a_241_164# 0.11fF
C252 g0 a_140_n252# 0.12fF
C253 g3 a_98_139# 0.25fF
C254 w_52_200# vdd 0.09fF
C255 w_163_225# g1 0.07fF
C256 w_n69_84# vdd 0.09fF
C257 a_241_164# a_145_231# 0.07fF
C258 p0 a_76_n182# 0.08fF
C259 w_166_68# vdd 0.09fF
C260 w_n65_145# p3 0.07fF
C261 g0 m1_163_n48# 0.02fF
C262 a_148_74# vdd 1.34fF
C263 w_n69_180# p3 0.07fF
C264 w_477_45# vdd 0.09fF
C265 a_426_70# a_472_117# 0.31fF
C266 a_106_n9# vdd 2.64fF
C267 a3 a_n266_193# 0.07fF
C268 a_42_58# gnd 0.03fF
C269 g1 a_177_137# 0.01fF
C270 a_98_139# a_542_198# 0.04fF
C271 w_n69_212# a_n133_157# 0.07fF
C272 w_n201_187# b3 0.07fF
C273 w_n201_155# a_n266_193# 0.07fF
C274 w_52_200# a_34_206# 0.07fF
C275 w_n201_27# g2 0.07fF
C276 w_n201_n69# vdd 0.09fF
C277 w_28_52# p2 0.07fF
C278 w_60_52# g1 0.07fF
C279 w_563_192# a_542_198# 0.25fF
C280 p3 a_298_139# 0.07fF
C281 c3 vdd 0.45fF
C282 g1 p1 0.68fF
C283 p2 g0 0.74fF
C284 w_316_133# g0 0.07fF
C285 w_729_113# p3 0.07fF
C286 a_140_n155# a_279_n316# 0.98fF
C287 w_131_225# p3 0.07fF
C288 c0 s0 0.95fF
C289 w_564_n242# c3 0.07fF
C290 a_459_51# vdd 2.23fF
C291 p0 a_653_n389# 0.08fF
C292 g1 a_42_58# 0.48fF
C293 w_630_183# c4 0.07fF
C294 w_671_n328# c0 0.07fF
C295 a_577_198# a_472_117# 2.20fF
C296 g2 a_244_7# 0.22fF
C297 w_694_n36# s2 0.07fF
C298 w_639_n328# p0 0.07fF
C299 a_140_n155# vdd 1.04fF
C300 a_n133_n99# gnd 0.47fF
C301 w_n69_52# a2 0.07fF
C302 w_166_68# g0 0.07fF
C303 w_62_n94# vdd 0.09fF
C304 g0 a_148_74# 0.37fF
C305 p3 c0 1.52fF
C306 a_n266_n183# gnd 0.69fF
C307 w_n69_n172# a_n133_n227# 0.07fF
C308 g0 a_106_n9# 0.05fF
C309 w_404_n55# vdd 0.09fF
C310 w_230_68# a_244_7# 0.07fF
C311 g2 a_418_n118# 0.00fF
C312 w_n201_n165# vdd 0.09fF
C313 a_148_74# a_148_n14# 0.19fF
C314 a_106_n9# a_148_n14# 0.25fF
C315 p1 p0 1.09fF
C316 w_n201_n37# a1 0.07fF
C317 g0 a_140_n155# 0.11fF
C318 p1 b1 0.95fF
C319 w_729_n32# p2 0.07fF
C320 a_322_n165# a_354_n165# 0.82fF
C321 w_573_45# a_459_51# 0.07fF
C322 w_30_n94# p1 0.07fF
C323 a_676_48# s3 1.05fF
C324 w_n69_n204# b0 0.07fF
C325 w_n201_n69# a_n266_n63# 0.07fF
C326 a1 b1 0.23fF
C327 c2 c1 0.34fF
C328 a_676_n97# s2 1.05fF
C329 w_265_n249# a_240_n171# 0.07fF
C330 c0 a_44_n88# 0.54fF
C331 a_240_n171# gnd 0.41fF
C332 a_n133_n99# b1 0.40fF
C333 a_459_n85# gnd 1.38fF
C334 w_367_n256# c2 0.07fF
C335 w_n69_n76# b1 0.07fF
C336 g1 a_240_n171# 0.04fF
C337 c1 gnd 0.41fF
C338 w_300_n249# a_279_n243# 0.11fF
C339 w_194_n110# c0 0.01fF
C340 p2 a_354_n165# 0.08fF
C341 w_462_n235# a_441_n229# 0.13fF
C342 w_195_n258# vdd 0.09fF
C343 w_639_n183# a_653_n244# 0.07fF
C344 p2 s2 0.55fF
C345 w_n201_n165# a0 0.07fF
C346 a_n266_n183# a_n266_n191# 0.42fF
C347 w_639_n328# a_653_n389# 0.07fF
C348 g1 a_314_n243# 0.05fF
C349 g0 a_176_n172# 0.07fF
C350 w_195_225# vdd 0.09fF
C351 p3 vdd 0.74fF
C352 p1 a_523_n91# 0.01fF
C353 a_241_164# gnd 0.51fF
C354 g3 a_426_70# 0.00fF
C355 g0 a_140_n320# 0.05fF
C356 g2 gnd 0.41fF
C357 w_227_225# a_241_164# 0.07fF
C358 w_n201_91# vdd 0.08fF
C359 c0 b0 0.08fF
C360 a_34_138# gnd 0.69fF
C361 a_472_198# vdd 2.13fF
C362 a_98_139# p3 0.63fF
C363 p0 a_240_n171# 0.06fF
C364 w_598_192# a_605_159# 0.07fF
C365 w_92_52# vdd 0.09fF
C366 a_298_139# vdd 1.79fF
C367 p0 a_459_n85# 0.01fF
C368 p2 a_145_231# 0.88fF
C369 g1 g2 0.51fF
C370 g3 b3 0.31fF
C371 c0 a_491_n91# 0.01fF
C372 a_472_117# gnd 2.31fF
C373 p3 a_34_206# 0.07fF
C374 a_241_164# a_507_198# 0.02fF
C375 p0 c1 0.05fF
C376 w_131_225# vdd 0.09fF
C377 a_244_7# a_441_n306# 0.31fF
C378 a_n133_29# vdd 0.96fF
C379 a_n266_73# gnd 0.69fF
C380 c0 a_44_n241# 0.48fF
C381 w_n201_187# a_n266_193# 0.07fF
C382 w_528_192# a_507_198# 0.25fF
C383 a_n133_157# b3 0.40fF
C384 p3 g0 0.00fF
C385 a_42_n10# gnd 0.69fF
C386 w_662_109# p3 0.07fF
C387 w_226_n110# a_240_n171# 0.07fF
C388 c0 vdd 0.38fF
C389 p2 a2 0.55fF
C390 w_n69_n204# a0 0.07fF
C391 w_607_45# a_605_159# 0.07fF
C392 w_412_133# a_298_139# 0.07fF
C393 g1 a_42_n10# 0.07fF
C394 a_44_n88# vdd 1.37fF
C395 w_335_n249# a_140_n155# 0.07fF
C396 p2 a_244_7# 0.95fF
C397 w_694_n36# c2 0.07fF
C398 a_507_198# a_472_117# 0.12fF
C399 a_542_198# a_577_198# 2.13fF
C400 w_662_n36# a_676_n97# 0.07fF
C401 a_418_n118# a_441_n306# 0.26fF
C402 a_n266_n55# gnd 0.69fF
C403 g2 b2 0.31fF
C404 w_n201_n101# g1 0.07fF
C405 w_n201_91# a_n266_65# 0.07fF
C406 w_n69_84# a2 0.07fF
C407 g0 a_298_139# 0.32fF
C408 a_98_139# c0 2.15fF
C409 a_472_117# c4 0.07fF
C410 a_176_n104# gnd 0.03fF
C411 w_198_68# a_148_74# 0.07fF
C412 w_60_52# a_42_58# 0.07fF
C413 w_n69_52# b2 0.07fF
C414 w_340_n55# vdd 0.09fF
C415 g2 p0 0.06fF
C416 p2 a_290_n49# 0.27fF
C417 a_148_74# a_244_7# 0.07fF
C418 g0 a_180_n20# 0.01fF
C419 w_194_n110# vdd 0.09fF
C420 p1 a1 0.55fF
C421 a_n266_73# b2 0.07fF
C422 a_106_n9# a_244_7# 0.30fF
C423 g0 c0 0.16fF
C424 p1 a_362_23# 0.01fF
C425 p1 a_n133_n99# 1.05fF
C426 a_148_n14# a_180_n20# 0.62fF
C427 w_662_n36# p2 0.07fF
C428 a_290_n159# a_322_n165# 0.82fF
C429 w_509_45# a_459_51# 0.07fF
C430 w_n69_n76# p1 0.07fF
C431 c3 a_676_48# 0.40fF
C432 a1 a_n133_n99# 0.08fF
C433 a_106_n9# a_418_n118# 0.29fF
C434 c2 a_676_n97# 0.40fF
C435 w_162_n110# p1 0.17fF
C436 w_194_n110# g0 0.07fF
C437 w_n69_n76# a1 0.07fF
C438 w_n201_n229# vdd 0.09fF
C439 a_n266_n55# b1 0.07fF
C440 w_94_n247# a_108_n308# 0.07fF
C441 a_44_n241# vdd 0.89fF
C442 a_676_n97# gnd 0.47fF
C443 w_404_n55# a_290_n49# 0.07fF
C444 w_126_n258# vdd 0.09fF
C445 a_511_n229# a_441_n306# 0.98fF
C446 w_404_n55# a_418_n118# 0.07fF
C447 a_441_n306# gnd 1.85fF
C448 p2 c2 0.81fF
C449 w_427_n235# vdd 0.13fF
C450 w_532_n235# a_441_n306# 0.11fF
C451 w_226_n110# a_176_n104# 0.07fF
C452 w_n201_n229# g0 0.07fF
C453 w_564_n242# vdd 0.09fF
C454 p1 a_240_n171# 0.28fF
C455 w_300_n249# g1 0.07fF
C456 a_98_139# vdd 2.12fF
C457 g3 gnd 0.41fF
C458 g2 a_441_n229# 0.01fF
C459 p1 c1 0.15fF
C460 a_34_206# vdd 0.89fF
C461 w_n69_212# vdd 0.09fF
C462 w_412_133# vdd 0.09fF
C463 a_426_70# p3 0.03fF
C464 w_126_n258# g0 0.20fF
C465 a_241_164# a_605_159# 0.03fF
C466 c0 a_44_n176# 0.10fF
C467 a_n133_157# gnd 0.47fF
C468 w_28_52# vdd 0.09fF
C469 w_563_192# a_98_139# 0.07fF
C470 w_195_225# a_145_231# 0.07fF
C471 g1 p2 0.15fF
C472 p1 s1 0.55fF
C473 a_44_n88# a_44_n176# 0.19fF
C474 g3 a_n266_193# 0.07fF
C475 a_98_139# a_34_206# 0.07fF
C476 g0 vdd 1.13fF
C477 p3 a_145_231# 0.07fF
C478 c3 c2 0.24fF
C479 w_n201_n197# a_n266_n191# 0.07fF
C480 w_662_109# vdd 0.09fF
C481 p3 b3 0.95fF
C482 a_426_70# a_472_198# 0.02fF
C483 a_244_7# a_476_n229# 0.05fF
C484 a_148_74# gnd 0.03fF
C485 w_706_n179# p1 0.07fF
C486 a_106_n9# a_511_n229# 0.05fF
C487 a_n266_65# vdd 0.89fF
C488 a0 b0 0.23fF
C489 w_n65_145# b3 0.07fF
C490 w_493_192# a_472_198# 0.25fF
C491 w_573_45# vdd 0.09fF
C492 w_62_n247# c0 0.07fF
C493 a_n266_201# b3 0.07fF
C494 a_605_159# a_472_117# 0.36fF
C495 a_426_70# a_298_139# 0.07fF
C496 a_106_n9# gnd 0.67fF
C497 w_30_n247# p0 0.18fF
C498 w_n69_180# b3 0.07fF
C499 w_598_192# a_472_117# 0.23fF
C500 w_134_68# p2 0.07fF
C501 g2 p1 0.28fF
C502 c3 gnd 0.41fF
C503 w_630_183# a_472_117# 0.07fF
C504 w_348_133# a_298_139# 0.07fF
C505 a_n266_n63# vdd 0.89fF
C506 a_459_51# gnd 0.45fF
C507 p2 b2 0.95fF
C508 g1 a_106_n9# 0.47fF
C509 a_507_198# a_542_198# 2.13fF
C510 w_131_225# a_145_231# 0.07fF
C511 w_n201_91# a2 0.07fF
C512 a_426_70# c0 0.07fF
C513 a_140_n155# gnd 1.05fF
C514 p3 a_676_48# 0.08fF
C515 w_134_68# a_148_74# 0.07fF
C516 p2 p0 0.37fF
C517 w_276_n55# vdd 0.09fF
C518 g0 a_148_n14# 0.10fF
C519 b3 c0 0.08fF
C520 g1 a_140_n155# 0.05fF
C521 a2 a_n133_29# 0.08fF
C522 w_n65_17# a2 0.07fF
C523 g0 a_330_23# 0.01fF
C524 a_42_58# a_42_n10# 0.42fF
C525 w_694_109# s3 0.07fF
C526 w_372_n55# p2 0.07fF
C527 w_445_45# a_459_51# 0.07fF
C528 a_106_n9# p0 0.08fF
C529 p1 a_176_n104# 0.07fF
C530 w_n201_n69# b1 0.07fF
C531 p0 a_459_51# 0.25fF
C532 c0 a_290_n49# 0.32fF
C533 a_44_n176# vdd 0.25fF
C534 p0 a_140_n155# 0.06fF
C535 a_176_n172# gnd 0.69fF
C536 w_62_n247# a_44_n241# 0.07fF
C537 a_108_n308# a_140_n252# 0.07fF
C538 w_94_n94# c0 0.01fF
C539 w_163_n258# a_140_n252# 0.09fF
C540 a_555_n91# gnd 0.25fF
C541 a_279_n243# a_279_n316# 0.12fF
C542 c1 s1 0.95fF
C543 w_94_n94# a_44_n88# 0.07fF
C544 w_340_n55# a_290_n49# 0.07fF
C545 a_476_n229# a_511_n229# 0.90fF
C546 a_279_n243# vdd 0.69fF
C547 a_441_n229# a_441_n306# 0.12fF
C548 a_140_n320# gnd 0.89fF
C549 w_62_n247# vdd 0.09fF
C550 w_335_n249# a_279_n316# 0.09fF
C551 w_706_n179# c1 0.07fF
C552 p2 a_523_n91# 0.08fF
C553 w_497_n235# a_511_n229# 0.11fF
C554 a_653_n244# vdd 0.45fF
C555 w_162_n110# a_176_n104# 0.07fF
C556 w_706_n179# s1 0.07fF
C557 a_426_70# vdd 0.45fF
C558 p1 a_322_n165# 0.10fF
C559 w_706_n324# s0 0.07fF
C560 a_145_231# vdd 1.34fF
C561 w_n201_219# vdd 0.08fF
C562 w_n201_n165# a_n266_n191# 0.07fF
C563 w_348_133# vdd 0.09fF
C564 a_n266_201# gnd 0.69fF
C565 a_426_70# a_98_139# 0.20fF
C566 g3 a_605_159# 0.02fF
C567 w_84_200# vdd 0.09fF
C568 w_528_192# a_241_164# 0.07fF
C569 w_n201_27# vdd 0.07fF
C570 p3 g1 0.00fF
C571 c0 a_290_n159# 0.10fF
C572 w_n201_155# g3 0.07fF
C573 w_284_133# p3 0.07fF
C574 w_198_68# vdd 0.09fF
C575 w_412_133# a_426_70# 0.07fF
C576 w_639_n183# p1 0.07fF
C577 a_176_n104# a_240_n171# 0.07fF
C578 g0 m5_167_n48# 0.06fF
C579 p0 a_555_n91# 0.08fF
C580 w_20_200# p3 0.07fF
C581 w_84_200# a_98_139# 0.07fF
C582 w_509_45# vdd 0.09fF
C583 a_241_164# a_472_117# 0.83fF
C584 a_145_231# a_145_143# 0.19fF
C585 c0 a_44_n309# 0.07fF
C586 a_98_139# a_577_198# 0.05fF
C587 a_244_7# vdd 0.45fF
C588 a_n133_29# gnd 0.47fF
C589 w_n69_n204# p0 0.07fF
C590 g2 a_34_138# 0.07fF
C591 a_n266_201# a_n266_193# 0.42fF
C592 p2 a_177_137# 0.08fF
C593 a3 a_n133_157# 0.08fF
C594 w_84_200# a_34_206# 0.07fF
C595 w_563_192# a_577_198# 0.23fF
C596 w_n69_n44# vdd 0.09fF
C597 a_676_48# vdd 0.45fF
C598 p2 p1 0.68fF
C599 w_445_45# p3 0.07fF
C600 w_284_133# a_298_139# 0.07fF
C601 p2 a_42_58# 0.07fF
C602 a_472_198# a_507_198# 2.13fF
C603 a_290_n49# vdd 1.79fF
C604 p0 s0 0.55fF
C605 w_671_n328# p0 0.07fF
C606 w_729_n32# s2 0.07fF
C607 a_44_n88# gnd 0.03fF
C608 a_418_n118# vdd 0.45fF
C609 w_706_n324# c0 0.07fF
C610 w_n201_27# a_n266_65# 0.07fF
C611 p1 a_148_74# 0.88fF
C612 p3 p0 0.00fF
C613 p2 a_362_23# 0.08fF
C614 w_94_n94# vdd 0.09fF
C615 a_605_159# a_459_51# 0.07fF
C616 g1 c0 0.19fF
C617 a_n133_n227# b0 0.40fF
C618 p1 a_106_n9# 1.78fF
C619 a2 a_n266_65# 0.07fF
C620 w_662_n36# vdd 0.09fF
C621 a_n133_29# b2 0.40fF
C622 a_42_58# a_106_n9# 0.07fF
C623 a_298_139# a_298_29# 0.08fF
C624 p1 c3 0.63fF
C625 w_662_109# a_676_48# 0.07fF
C626 w_694_109# c3 0.07fF
C627 w_n65_17# b2 0.07fF
C628 p1 a_459_51# 0.73fF
C629 b2 c0 0.08fF
C630 p1 a_140_n155# 0.12fF
C631 a_n133_n227# vdd 0.96fF
C632 w_607_45# a_459_51# 0.07fF
C633 a_523_n91# a_555_n91# 1.03fF
C634 w_n65_n239# b0 0.07fF
C635 c0 p0 0.47fF
C636 a_322_n165# a_314_n243# 0.13fF
C637 p0 a_44_n88# 0.88fF
C638 c0 b1 0.08fF
C639 c2 a_279_n316# 0.07fF
C640 a_44_n241# a_44_n309# 0.42fF
C641 w_30_n94# c0 0.01fF
C642 w_163_n258# a_140_n320# 0.07fF
C643 c2 vdd 0.45fF
C644 a_491_n91# gnd 0.25fF
C645 w_276_n55# a_290_n49# 0.07fF
C646 w_30_n94# a_44_n88# 0.07fF
C647 w_n65_n111# b1 0.07fF
C648 w_300_n249# a_314_n243# 0.09fF
C649 a_441_n229# a_476_n229# 0.90fF
C650 a_44_n241# gnd 0.03fF
C651 w_226_n110# c0 0.01fF
C652 w_462_n235# a_476_n229# 0.11fF
C653 w_265_n249# vdd 0.11fF
C654 a_279_n316# gnd 1.42fF
C655 a_653_n389# s0 1.05fF
C656 vdd gnd 1.04fF
C657 g1 a_279_n316# 0.39fF
C658 w_227_225# vdd 0.09fF
C659 a_98_139# gnd 0.48fF
C660 g1 vdd 0.45fF
C661 w_284_133# vdd 0.09fF
C662 a0 a_n133_n227# 0.08fF
C663 g3 a_241_164# 0.00fF
C664 a_34_206# gnd 0.03fF
C665 a_n266_193# vdd 0.89fF
C666 w_20_200# vdd 0.09fF
C667 w_493_192# a_426_70# 0.07fF
C668 w_n201_59# vdd 0.09fF
C669 a_145_143# gnd 0.72fF
C670 a_605_159# p3 0.75fF
C671 c0 a_76_n182# 0.01fF
C672 p0 b0 0.95fF
C673 w_134_68# vdd 0.09fF
C674 c4 vdd 0.45fF
C675 c3 c1 0.16fF
C676 p2 g2 3.25fF
C677 a_140_n155# a_240_n171# 0.00fF
C678 g0 gnd 0.41fF
C679 p3 a3 0.55fF
C680 a_44_n88# a_76_n182# 0.62fF
C681 a_290_n49# a_354_n165# 0.82fF
C682 w_445_45# vdd 0.09fF
C683 w_n65_145# a3 0.07fF
C684 w_380_133# p2 0.07fF
C685 g1 a_145_143# 0.10fF
C686 a_241_164# a_542_198# 0.05fF
C687 a_n266_65# gnd 0.03fF
C688 p0 a_44_n241# 0.07fF
C689 w_52_200# g2 0.07fF
C690 w_20_200# a_34_206# 0.07fF
C691 w_n69_180# a3 0.07fF
C692 w_n69_52# p2 0.07fF
C693 w_528_192# a_542_198# 0.23fF
C694 w_n201_n37# vdd 0.09fF
C695 p3 p1 0.01fF
C696 a_148_n14# gnd 0.72fF
C697 g1 g0 0.35fF
C698 w_694_109# p3 0.07fF
C699 c0 a_653_n389# 0.39fF
C700 a_140_n155# a_314_n243# 0.02fF
C701 w_n65_n239# a0 0.07fF
C702 p0 vdd 0.03fF
C703 w_n201_n229# a_n266_n191# 0.07fF
C704 a_n266_n191# b0 0.48fF
C705 w_541_45# p2 0.07fF
C706 a_542_198# a_472_117# 0.12fF
C707 g2 a_106_n9# 0.07fF
C708 w_729_n32# c2 0.07fF
C709 a_n266_n63# gnd 0.03fF
C710 m5_167_n48# Gnd 0.03fF **FLOATING
C711 m1_163_n48# Gnd 0.02fF **FLOATING
C712 gnd Gnd 8.59fF
C713 s0 Gnd 0.36fF
C714 a_653_n389# Gnd 0.88fF
C715 vdd Gnd 5.32fF
C716 s1 Gnd 0.36fF
C717 a_653_n244# Gnd 0.88fF
C718 a_441_n306# Gnd 1.05fF
C719 a_511_n229# Gnd 0.42fF
C720 a_476_n229# Gnd 0.42fF
C721 a_441_n229# Gnd 0.42fF
C722 a_279_n316# Gnd 0.78fF
C723 a_314_n243# Gnd 0.36fF
C724 a_279_n243# Gnd 0.36fF
C725 a_140_n252# Gnd 0.35fF
C726 a_44_n309# Gnd 0.33fF
C727 a_140_n320# Gnd 1.07fF
C728 a_108_n308# Gnd 0.39fF
C729 a_44_n241# Gnd 0.54fF
C730 c1 Gnd 1.36fF
C731 s2 Gnd 0.36fF
C732 a_676_n97# Gnd 0.88fF
C733 c2 Gnd 1.38fF
C734 a_555_n91# Gnd 0.64fF
C735 a_523_n91# Gnd 0.64fF
C736 a_491_n91# Gnd 0.64fF
C737 a_459_n85# Gnd 0.65fF
C738 a_354_n165# Gnd 0.53fF
C739 a_322_n165# Gnd 0.53fF
C740 a_290_n159# Gnd 0.55fF
C741 a_176_n172# Gnd 0.02fF
C742 a_76_n182# Gnd 0.43fF
C743 b0 Gnd 1.25fF
C744 a_240_n171# Gnd 0.85fF
C745 a_44_n176# Gnd 0.45fF
C746 a_n133_n227# Gnd 0.88fF
C747 a_n266_n191# Gnd 0.54fF
C748 a_n266_n183# Gnd 0.33fF
C749 a0 Gnd 5.52fF
C750 a_176_n104# Gnd 0.54fF
C751 a_418_n118# Gnd 1.35fF
C752 a_140_n155# Gnd 2.92fF
C753 b1 Gnd 1.25fF
C754 a_44_n88# Gnd 0.69fF
C755 a_n133_n99# Gnd 0.88fF
C756 a_n266_n63# Gnd 0.54fF
C757 a_n266_n55# Gnd 0.33fF
C758 a_290_n49# Gnd 0.86fF
C759 a_459_51# Gnd 1.07fF
C760 p0 Gnd 10.58fF
C761 c0 Gnd 4.14fF
C762 a_362_23# Gnd 0.53fF
C763 a_330_23# Gnd 0.53fF
C764 s3 Gnd 0.36fF
C765 a_676_48# Gnd 0.88fF
C766 c3 Gnd 1.23fF
C767 a_298_29# Gnd 0.55fF
C768 a_180_n20# Gnd 0.43fF
C769 a1 Gnd 5.52fF
C770 a_148_n14# Gnd 0.45fF
C771 a_42_n10# Gnd 0.33fF
C772 a_244_7# Gnd 1.11fF
C773 a_106_n9# Gnd 5.39fF
C774 b2 Gnd 1.25fF
C775 a_n133_29# Gnd 0.88fF
C776 a_42_58# Gnd 0.54fF
C777 a_n266_65# Gnd 0.54fF
C778 a_n266_73# Gnd 0.33fF
C779 a2 Gnd 5.52fF
C780 a_148_74# Gnd 0.69fF
C781 c4 Gnd 0.38fF
C782 a_298_139# Gnd 0.86fF
C783 p1 Gnd 18.63fF
C784 g0 Gnd 7.33fF
C785 a_472_117# Gnd 1.34fF
C786 a_577_198# Gnd 0.77fF
C787 a_542_198# Gnd 0.77fF
C788 a_507_198# Gnd 0.77fF
C789 a_472_198# Gnd 0.77fF
C790 a_177_137# Gnd 0.43fF
C791 a_145_143# Gnd 0.45fF
C792 a_34_138# Gnd 0.33fF
C793 b3 Gnd 1.25fF
C794 a_n133_157# Gnd 0.88fF
C795 a_n266_193# Gnd 0.54fF
C796 a_n266_201# Gnd 0.33fF
C797 a3 Gnd 5.52fF
C798 a_34_206# Gnd 0.54fF
C799 g2 Gnd 8.48fF
C800 a_145_231# Gnd 0.69fF
C801 p2 Gnd 15.33fF
C802 g1 Gnd 7.22fF
C803 p3 Gnd 8.53fF
C804 a_605_159# Gnd 2.15fF
C805 a_98_139# Gnd 2.34fF
C806 a_241_164# Gnd 1.83fF
C807 a_426_70# Gnd 0.72fF
C808 g3 Gnd 6.69fF
C809 w_706_n324# Gnd 1.36fF
C810 w_671_n328# Gnd 1.36fF
C811 w_639_n328# Gnd 1.36fF
C812 w_564_n242# Gnd 1.36fF
C813 w_706_n179# Gnd 1.36fF
C814 w_671_n183# Gnd 1.36fF
C815 w_639_n183# Gnd 1.36fF
C816 w_532_n235# Gnd 2.40fF
C817 w_497_n235# Gnd 2.40fF
C818 w_462_n235# Gnd 2.40fF
C819 w_427_n235# Gnd 2.40fF
C820 w_367_n256# Gnd 1.36fF
C821 w_335_n249# Gnd 1.88fF
C822 w_300_n249# Gnd 1.88fF
C823 w_265_n249# Gnd 1.88fF
C824 w_195_n258# Gnd 1.36fF
C825 w_163_n258# Gnd 1.36fF
C826 w_126_n258# Gnd 1.36fF
C827 w_94_n247# Gnd 1.36fF
C828 w_62_n247# Gnd 1.36fF
C829 w_30_n247# Gnd 1.36fF
C830 w_n65_n239# Gnd 1.36fF
C831 w_n69_n204# Gnd 1.36fF
C832 w_n201_n229# Gnd 1.36fF
C833 w_n69_n172# Gnd 1.36fF
C834 w_n201_n197# Gnd 1.36fF
C835 w_n201_n165# Gnd 1.36fF
C836 w_226_n110# Gnd 1.36fF
C837 w_194_n110# Gnd 1.36fF
C838 w_162_n110# Gnd 1.36fF
C839 w_729_n32# Gnd 1.36fF
C840 w_694_n36# Gnd 1.36fF
C841 w_662_n36# Gnd 1.36fF
C842 w_404_n55# Gnd 1.36fF
C843 w_372_n55# Gnd 1.36fF
C844 w_340_n55# Gnd 1.36fF
C845 w_308_n55# Gnd 1.36fF
C846 w_276_n55# Gnd 1.36fF
C847 w_126_n94# Gnd 1.36fF
C848 w_94_n94# Gnd 1.36fF
C849 w_62_n94# Gnd 1.36fF
C850 w_30_n94# Gnd 1.36fF
C851 w_n65_n111# Gnd 1.36fF
C852 w_n69_n76# Gnd 1.36fF
C853 w_n201_n101# Gnd 1.36fF
C854 w_n69_n44# Gnd 1.36fF
C855 w_n201_n69# Gnd 1.36fF
C856 w_n201_n37# Gnd 1.36fF
C857 w_n65_17# Gnd 1.36fF
C858 w_607_45# Gnd 1.36fF
C859 w_573_45# Gnd 1.36fF
C860 w_541_45# Gnd 1.36fF
C861 w_509_45# Gnd 1.36fF
C862 w_477_45# Gnd 1.36fF
C863 w_445_45# Gnd 1.36fF
C864 w_729_113# Gnd 1.36fF
C865 w_694_109# Gnd 1.36fF
C866 w_662_109# Gnd 1.36fF
C867 w_230_68# Gnd 1.36fF
C868 w_198_68# Gnd 1.36fF
C869 w_166_68# Gnd 1.36fF
C870 w_134_68# Gnd 1.36fF
C871 w_92_52# Gnd 1.36fF
C872 w_60_52# Gnd 1.36fF
C873 w_28_52# Gnd 1.36fF
C874 w_n69_52# Gnd 1.36fF
C875 w_n201_27# Gnd 1.36fF
C876 w_n69_84# Gnd 1.36fF
C877 w_n201_59# Gnd 1.36fF
C878 w_n201_91# Gnd 1.36fF
C879 w_630_183# Gnd 1.36fF
C880 w_412_133# Gnd 1.36fF
C881 w_380_133# Gnd 1.36fF
C882 w_348_133# Gnd 1.36fF
C883 w_316_133# Gnd 1.36fF
C884 w_284_133# Gnd 1.36fF
C885 w_n65_145# Gnd 1.36fF
C886 w_598_192# Gnd 5.51fF
C887 w_563_192# Gnd 5.51fF
C888 w_528_192# Gnd 5.51fF
C889 w_493_192# Gnd 5.51fF
C890 w_458_192# Gnd 5.51fF
C891 w_227_225# Gnd 1.36fF
C892 w_195_225# Gnd 1.36fF
C893 w_163_225# Gnd 1.36fF
C894 w_131_225# Gnd 1.36fF
C895 w_84_200# Gnd 1.36fF
C896 w_52_200# Gnd 1.36fF
C897 w_20_200# Gnd 1.36fF
C898 w_n69_180# Gnd 1.36fF
C899 w_n201_155# Gnd 1.36fF
C900 w_n69_212# Gnd 1.36fF
C901 w_n201_187# Gnd 1.36fF
C902 w_n201_219# Gnd 1.36fF
