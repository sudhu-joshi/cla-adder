.include TSMC_180nm.txt
.include subckt.txt

.param SUPPLY=1.8
.param LAMBDA = 0.09u
.param len = 2*LAMBDA
.param W_P = 20*LAMBDA
.param W_N = 10*LAMBDA

.global gnd vdd 
vdd vdd gnd 'SUPPLY'

* Input Pulses
VA A gnd pulse (0 SUPPLY 10ns .1ns .1ns 10ns 20ns)
VB B gnd pulse (0 SUPPLY 20ns .1ns .1ns 20ns 40ns)
VC C gnd pulse (0 SUPPLY 40ns .1ns .1ns 40ns 80ns)
VD D gnd pulse (0 SUPPLY 80ns .1ns .1ns 80ns 160ns)
Vclk clk gnd pulse (0 SUPPLY 5ns .1ns .1ns 5ns 10ns)

* .subckt d_latch q d en vdd gnd 
* * d_ff pos edge
.subckt d_block_4bit q3 q2 q1 q0 d3 d2 d1 d0 clk vdd gnd

Xd3_ff q3 d3 clk vdd gnd d_ff
Xd2_ff q2 d2 clk vdd gnd d_ff
Xd1_ff q1 d1 clk vdd gnd d_ff
Xd0_ff q0 d0 clk vdd gnd d_ff

.ends d_block_4bit


Xd_block_4bit out A clk vdd gnd d_block_4bit

* Simulation Setup
.tran 0.01ns 320ns
.control
    set hcopypscolor = 1
    set color0 = black
    set color1 = white
    run
    set curplottitle= d_block_4bit
    plot v(A) v(clk) v(out)+2

.endc
.end
