magic
tech scmos
timestamp 1732037632
<< nwell >>
rect -1 30 25 122
rect 34 30 60 122
rect 69 30 95 122
rect 104 30 130 122
rect 136 23 162 75
<< ntransistor >>
rect 11 -41 13 -1
rect 46 -42 48 -2
rect 81 -42 83 -2
rect 116 -42 118 -2
rect 148 -42 150 -2
<< ptransistor >>
rect 11 36 13 116
rect 46 36 48 116
rect 81 36 83 116
rect 116 36 118 116
rect 148 29 150 69
<< ndiffusion >>
rect 10 -41 11 -1
rect 13 -41 14 -1
rect 45 -42 46 -2
rect 48 -42 49 -2
rect 80 -42 81 -2
rect 83 -42 84 -2
rect 115 -42 116 -2
rect 118 -42 119 -2
rect 147 -42 148 -2
rect 150 -42 151 -2
<< pdiffusion >>
rect 10 36 11 116
rect 13 36 14 116
rect 45 36 46 116
rect 48 36 49 116
rect 80 36 81 116
rect 83 36 84 116
rect 115 36 116 116
rect 118 36 119 116
rect 147 29 148 69
rect 150 29 151 69
<< ndcontact >>
rect 5 -41 10 -1
rect 14 -41 19 -1
rect 40 -42 45 -2
rect 49 -42 54 -2
rect 75 -42 80 -2
rect 84 -42 89 -2
rect 110 -42 115 -2
rect 119 -42 124 -2
rect 142 -42 147 -2
rect 151 -42 156 -2
<< pdcontact >>
rect 5 36 10 116
rect 14 36 19 116
rect 40 36 45 116
rect 49 36 54 116
rect 75 36 80 116
rect 84 36 89 116
rect 110 36 115 116
rect 119 36 124 116
rect 142 29 147 69
rect 151 29 156 69
<< polysilicon >>
rect 11 116 13 120
rect 46 116 48 120
rect 81 116 83 120
rect 116 116 118 120
rect 148 69 150 73
rect 11 -1 13 36
rect 46 22 48 36
rect 81 22 83 36
rect 116 22 118 36
rect 46 -2 48 6
rect 81 -2 83 6
rect 116 -2 118 6
rect 148 -2 150 29
rect 11 -44 13 -41
rect 46 -45 48 -42
rect 81 -45 83 -42
rect 116 -45 118 -42
rect 148 -45 150 -42
<< polycontact >>
rect 6 19 11 24
rect 41 22 46 27
rect 76 22 81 27
rect 111 22 116 27
rect 143 13 148 18
rect 41 1 46 6
rect 76 1 81 6
rect 111 1 116 6
<< metal1 >>
rect -1 122 25 125
rect 28 122 60 125
rect 63 122 95 125
rect 98 122 130 125
rect 5 116 10 122
rect 14 26 19 36
rect 28 26 31 122
rect 40 116 45 122
rect -1 19 6 24
rect 14 23 31 26
rect 38 22 41 27
rect 49 26 54 36
rect 63 26 66 122
rect 75 116 80 122
rect 49 23 66 26
rect 73 22 76 27
rect 84 26 89 36
rect 98 26 101 122
rect 110 116 115 122
rect 136 75 162 78
rect 84 23 101 26
rect 105 22 111 27
rect 119 18 124 36
rect 142 69 147 75
rect 119 17 143 18
rect 14 14 143 17
rect 14 -1 19 14
rect 38 1 41 6
rect 49 -2 54 14
rect 73 1 76 6
rect 84 -2 89 14
rect 119 13 143 14
rect 151 15 156 29
rect 105 1 111 6
rect 119 -2 124 13
rect 151 10 162 15
rect 151 -2 156 10
rect 5 -46 10 -41
rect 40 -46 45 -42
rect 75 -46 80 -42
rect 110 -46 115 -42
rect 142 -46 147 -42
rect 5 -49 147 -46
<< metal2 >>
rect 70 14 73 27
rect -1 11 73 14
rect 70 1 73 11
<< metal3 >>
rect 35 18 38 27
rect -1 15 38 18
rect 35 1 38 15
<< metal4 >>
rect 105 10 108 27
rect -1 7 108 10
rect 105 1 108 7
<< pad >>
rect 35 22 41 27
rect 70 22 76 27
rect 105 22 111 27
rect 35 1 41 6
rect 70 1 76 6
rect 105 1 111 6
<< labels >>
rlabel metal1 -1 19 6 24 3 a
rlabel metal1 151 2 156 29 1 out
rlabel metal1 136 75 162 78 1 vdd!
rlabel metal1 5 -49 147 -46 1 gnd!
rlabel metal3 -1 15 38 18 1 b
rlabel metal2 -1 11 73 14 1 c
rlabel metal4 -1 7 108 10 1 d
rlabel metal1 -1 122 25 125 5 vdd!
<< end >>
