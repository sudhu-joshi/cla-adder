.include TSMC_180nm.txt
.include subckt.txt

.param SUPPLY=1.8
.param LAMBDA = 0.09u
.param len = 2*LAMBDA
.param W_P = 20*LAMBDA
.param W_N = 10*LAMBDA

.global gnd vdd 
vdd vdd gnd 'SUPPLY'

* Input Pulses
VA A gnd pulse (0 SUPPLY 10ns .1ns .1ns 10ns 20ns)
VB B gnd pulse (0 SUPPLY 20ns .1ns .1ns 20ns 40ns)
VC C gnd pulse (0 SUPPLY 40ns .1ns .1ns 40ns 80ns)
* VD D gnd pulse (0 SUPPLY 80ns .1ns .1ns 80ns 160ns)

* SPICE3 file created from and3.ext - technology: scmos

.option scale=0.09u

M1000 a_13_n32# a gnd gnd CMOSN w=40 l=2
+  ad=480 pd=184 as=480 ps=184
M1001 a_13_36# b vdd w_31_30# CMOSP w=40 l=2
+  ad=720 pd=276 as=960 ps=368
M1002 out a_13_36# vdd w_95_30# CMOSP w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1003 out a_13_36# gnd gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1004 a_13_36# c a_45_n38# gnd CMOSN w=40 l=2
+  ad=240 pd=92 as=480 ps=184
M1005 a_13_36# a vdd w_n1_30# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_13_36# c vdd w_63_30# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_45_n38# b a_13_n32# gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
C0 b c 0.05fF
C1 a a_13_36# 0.07fF
C2 w_95_30# vdd 0.09fF
C3 w_31_30# a_13_36# 0.07fF
C4 w_n1_30# vdd 0.09fF
C5 w_63_30# c 0.07fF
C6 a_13_n32# gnd 0.51fF
C7 a_13_36# gnd 0.03fF
C8 a_13_36# out 0.07fF
C9 b a_45_n38# 0.01fF
C10 c a_13_36# 0.85fF
C11 w_63_30# vdd 0.09fF
C12 a c 0.00fF
C13 w_95_30# a_13_36# 0.07fF
C14 w_n1_30# a_13_36# 0.07fF
C15 w_n1_30# a 0.07fF
C16 out gnd 0.44fF
C17 a_13_n32# a_45_n38# 0.41fF
C18 a_13_36# a_45_n38# 0.41fF
C19 a_13_36# vdd 1.34fF
C20 b a_13_n32# 0.10fF
C21 b a_13_36# 0.35fF
C22 w_95_30# out 0.07fF
C23 w_63_30# a_13_36# 0.07fF
C24 w_31_30# vdd 0.09fF
C25 a b 0.00fF
C26 w_31_30# b 0.07fF
C27 c a_45_n38# 0.10fF
C28 a_13_36# a_13_n32# 0.19fF
C29 vdd out 0.45fF
C30 gnd gnd 0.24fF
C31 a_45_n38# gnd 0.25fF
C32 a_13_n32# gnd 0.34fF
C33 out gnd 0.13fF
C34 vdd gnd 0.26fF
C35 a_13_36# gnd 0.67fF
C36 c gnd 1.00fF
C37 b gnd 0.38fF
C38 a gnd 0.23fF
C39 w_95_30# gnd 1.36fF
C40 w_63_30# gnd 1.36fF
C41 w_31_30# gnd 1.36fF
C42 w_n1_30# gnd 1.36fF


* Simulation Setup
.tran 0.01ns 170ns
.control
    set hcopypscolor = 1
    set color0 = black
    set color1 = white
    run
    set curplottitle= and3_post
    plot v(A) v(B)+2 v(C)+4 v(out)+6

.endc
.end



